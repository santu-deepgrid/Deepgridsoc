module dpram_be_256_256_8_8_128_128
  (input  [7:0] address_a,
   input  [15:0] byteena_a,
   input  clock0,
   input  [127:0] data_a,
   input  wren_a,
   input  [7:0] address_b,
   output [127:0] q_b);
  wire [127:0] q;
  wire [127:0] data;
  wire [7:0] address_r;
  wire [7:0] n45279_o;
  wire [7:0] n45280_o;
  wire [7:0] n45281_o;
  wire [7:0] n45282_o;
  wire [7:0] n45283_o;
  wire [7:0] n45284_o;
  wire [7:0] n45285_o;
  wire [7:0] n45286_o;
  wire [7:0] n45287_o;
  wire [7:0] n45288_o;
  wire [7:0] n45289_o;
  wire [7:0] n45290_o;
  wire [7:0] n45291_o;
  wire [7:0] n45292_o;
  wire [7:0] n45293_o;
  wire [7:0] n45294_o;
  wire [7:0] n45295_o;
  wire [7:0] n45296_o;
  wire [7:0] n45297_o;
  wire [7:0] n45298_o;
  wire [7:0] n45299_o;
  wire [7:0] n45300_o;
  wire [7:0] n45301_o;
  wire [7:0] n45302_o;
  wire [7:0] n45303_o;
  wire [7:0] n45304_o;
  wire [7:0] n45305_o;
  wire [7:0] n45306_o;
  wire [7:0] n45307_o;
  wire [7:0] n45308_o;
  wire [7:0] n45309_o;
  wire [7:0] n45310_o;
  wire n45314_o;
  wire [7:0] n45319_o;
  wire n45322_o;
  wire [7:0] n45327_o;
  wire n45330_o;
  wire [7:0] n45335_o;
  wire n45338_o;
  wire [7:0] n45343_o;
  wire n45346_o;
  wire [7:0] n45351_o;
  wire n45354_o;
  wire [7:0] n45359_o;
  wire n45362_o;
  wire [7:0] n45367_o;
  wire n45370_o;
  wire [7:0] n45375_o;
  wire n45378_o;
  wire [7:0] n45383_o;
  wire n45386_o;
  wire [7:0] n45391_o;
  wire n45394_o;
  wire [7:0] n45399_o;
  wire n45402_o;
  wire [7:0] n45407_o;
  wire n45410_o;
  wire [7:0] n45415_o;
  wire n45418_o;
  wire [7:0] n45423_o;
  wire n45426_o;
  wire [7:0] n45431_o;
  wire n45434_o;
  wire [7:0] n45439_o;
  wire n45446_o;
  wire n45448_o;
  wire n45450_o;
  wire n45452_o;
  wire n45454_o;
  wire n45456_o;
  wire n45458_o;
  wire n45460_o;
  wire n45462_o;
  wire n45464_o;
  wire n45466_o;
  wire n45468_o;
  wire n45470_o;
  wire n45472_o;
  wire n45474_o;
  wire n45476_o;
  wire [127:0] n45479_o;
  reg [7:0] n45480_q;
  wire [127:0] n45481_o;
  wire [7:0] n45482_data; // mem_rd
  wire [7:0] n45483_data; // mem_rd
  wire [7:0] n45484_data; // mem_rd
  wire [7:0] n45485_data; // mem_rd
  wire [7:0] n45486_data; // mem_rd
  wire [7:0] n45487_data; // mem_rd
  wire [7:0] n45488_data; // mem_rd
  wire [7:0] n45489_data; // mem_rd
  wire [7:0] n45490_data; // mem_rd
  wire [7:0] n45491_data; // mem_rd
  wire [7:0] n45492_data; // mem_rd
  wire [7:0] n45493_data; // mem_rd
  wire [7:0] n45494_data; // mem_rd
  wire [7:0] n45495_data; // mem_rd
  wire [7:0] n45496_data; // mem_rd
  wire [7:0] n45497_data; // mem_rd
  wire [127:0] n45498_o;
  assign q_b = n45481_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:55:8  */
  assign q = n45498_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:56:8  */
  assign data = n45479_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:57:8  */
  assign address_r = n45480_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45279_o = q[127:120];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45280_o = q[119:112];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45281_o = q[111:104];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45282_o = q[103:96];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45283_o = q[95:88];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45284_o = q[87:80];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45285_o = q[79:72];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45286_o = q[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45287_o = q[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45288_o = q[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45289_o = q[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45290_o = q[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45291_o = q[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45292_o = q[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45293_o = q[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45294_o = q[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45295_o = data_a[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45296_o = data_a[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45297_o = data_a[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45298_o = data_a[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45299_o = data_a[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45300_o = data_a[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45301_o = data_a[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45302_o = data_a[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45303_o = data_a[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45304_o = data_a[79:72];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45305_o = data_a[87:80];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45306_o = data_a[95:88];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45307_o = data_a[103:96];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45308_o = data_a[111:104];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45309_o = data_a[119:112];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45310_o = data_a[127:120];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45314_o = byteena_a[0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45319_o = data[127:120];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45322_o = byteena_a[1];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45327_o = data[119:112];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45330_o = byteena_a[2];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45335_o = data[111:104];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45338_o = byteena_a[3];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45343_o = data[103:96];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45346_o = byteena_a[4];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45351_o = data[95:88];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45354_o = byteena_a[5];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45359_o = data[87:80];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45362_o = byteena_a[6];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45367_o = data[79:72];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45370_o = byteena_a[7];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45375_o = data[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45378_o = byteena_a[8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45383_o = data[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45386_o = byteena_a[9];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45391_o = data[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45394_o = byteena_a[10];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45399_o = data[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45402_o = byteena_a[11];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45407_o = data[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45410_o = byteena_a[12];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45415_o = data[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45418_o = byteena_a[13];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45423_o = data[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45426_o = byteena_a[14];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45431_o = data[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45434_o = byteena_a[15];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45439_o = data[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45446_o = wren_a & n45434_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45448_o = wren_a & n45426_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45450_o = wren_a & n45418_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45452_o = wren_a & n45410_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45454_o = wren_a & n45402_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45456_o = wren_a & n45394_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45458_o = wren_a & n45386_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45460_o = wren_a & n45378_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45462_o = wren_a & n45370_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45464_o = wren_a & n45362_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45466_o = wren_a & n45354_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45468_o = wren_a & n45346_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45470_o = wren_a & n45338_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45472_o = wren_a & n45330_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45474_o = wren_a & n45322_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45476_o = wren_a & n45314_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n45479_o = {n45295_o, n45296_o, n45297_o, n45298_o, n45299_o, n45300_o, n45301_o, n45302_o, n45303_o, n45304_o, n45305_o, n45306_o, n45307_o, n45308_o, n45309_o, n45310_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  always @(posedge clock0)
    n45480_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n45481_o = {n45294_o, n45293_o, n45292_o, n45291_o, n45290_o, n45289_o, n45288_o, n45287_o, n45286_o, n45285_o, n45284_o, n45283_o, n45282_o, n45281_o, n45280_o, n45279_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n1[255:0] ; // memory
  assign n45482_data = ram_block_n1[address_r];
  always @(posedge clock0)
    if (n45446_o)
      ram_block_n1[address_a] <= n45439_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n2[255:0] ; // memory
  assign n45483_data = ram_block_n2[address_r];
  always @(posedge clock0)
    if (n45448_o)
      ram_block_n2[address_a] <= n45431_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n3[255:0] ; // memory
  assign n45484_data = ram_block_n3[address_r];
  always @(posedge clock0)
    if (n45450_o)
      ram_block_n3[address_a] <= n45423_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n4[255:0] ; // memory
  assign n45485_data = ram_block_n4[address_r];
  always @(posedge clock0)
    if (n45452_o)
      ram_block_n4[address_a] <= n45415_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n5[255:0] ; // memory
  assign n45486_data = ram_block_n5[address_r];
  always @(posedge clock0)
    if (n45454_o)
      ram_block_n5[address_a] <= n45407_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n6[255:0] ; // memory
  assign n45487_data = ram_block_n6[address_r];
  always @(posedge clock0)
    if (n45456_o)
      ram_block_n6[address_a] <= n45399_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n7[255:0] ; // memory
  assign n45488_data = ram_block_n7[address_r];
  always @(posedge clock0)
    if (n45458_o)
      ram_block_n7[address_a] <= n45391_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n8[255:0] ; // memory
  assign n45489_data = ram_block_n8[address_r];
  always @(posedge clock0)
    if (n45460_o)
      ram_block_n8[address_a] <= n45383_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n9[255:0] ; // memory
  assign n45490_data = ram_block_n9[address_r];
  always @(posedge clock0)
    if (n45462_o)
      ram_block_n9[address_a] <= n45375_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n10[255:0] ; // memory
  assign n45491_data = ram_block_n10[address_r];
  always @(posedge clock0)
    if (n45464_o)
      ram_block_n10[address_a] <= n45367_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n11[255:0] ; // memory
  assign n45492_data = ram_block_n11[address_r];
  always @(posedge clock0)
    if (n45466_o)
      ram_block_n11[address_a] <= n45359_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n12[255:0] ; // memory
  assign n45493_data = ram_block_n12[address_r];
  always @(posedge clock0)
    if (n45468_o)
      ram_block_n12[address_a] <= n45351_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n13[255:0] ; // memory
  assign n45494_data = ram_block_n13[address_r];
  always @(posedge clock0)
    if (n45470_o)
      ram_block_n13[address_a] <= n45343_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n14[255:0] ; // memory
  assign n45495_data = ram_block_n14[address_r];
  always @(posedge clock0)
    if (n45472_o)
      ram_block_n14[address_a] <= n45335_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n15[255:0] ; // memory
  assign n45496_data = ram_block_n15[address_r];
  always @(posedge clock0)
    if (n45474_o)
      ram_block_n15[address_a] <= n45327_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n16[255:0] ; // memory
  assign n45497_data = ram_block_n16[address_r];
  always @(posedge clock0)
    if (n45476_o)
      ram_block_n16[address_a] <= n45319_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  assign n45498_o = {n45497_data, n45496_data, n45495_data, n45494_data, n45493_data, n45492_data, n45491_data, n45490_data, n45489_data, n45488_data, n45487_data, n45486_data, n45485_data, n45484_data, n45483_data, n45482_data};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
endmodule

module sync_latch_128
  (input  enable_in,
   input  [127:0] data_in,
   output [127:0] data_out);
  wire [127:0] data_r;
  wire [127:0] n45271_o;
  assign data_out = data_r;
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:39:10  */
  assign data_r = n45271_o; // (signal)
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:45:4  */
  assign n45271_o = enable_in ? data_in : 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endmodule

module dpram_be_64_64_6_6_72_72
  (input  [5:0] address_a,
   input  [8:0] byteena_a,
   input  clock0,
   input  [71:0] data_a,
   input  wren_a,
   input  [5:0] address_b,
   output [71:0] q_b);
  wire [71:0] q;
  wire [71:0] data;
  wire [5:0] address_r;
  wire [7:0] n45129_o;
  wire [7:0] n45130_o;
  wire [7:0] n45131_o;
  wire [7:0] n45132_o;
  wire [7:0] n45133_o;
  wire [7:0] n45134_o;
  wire [7:0] n45135_o;
  wire [7:0] n45136_o;
  wire [7:0] n45137_o;
  wire [7:0] n45138_o;
  wire [7:0] n45139_o;
  wire [7:0] n45140_o;
  wire [7:0] n45141_o;
  wire [7:0] n45142_o;
  wire [7:0] n45143_o;
  wire [7:0] n45144_o;
  wire [7:0] n45145_o;
  wire [7:0] n45146_o;
  wire n45150_o;
  wire [7:0] n45155_o;
  wire n45158_o;
  wire [7:0] n45163_o;
  wire n45166_o;
  wire [7:0] n45171_o;
  wire n45174_o;
  wire [7:0] n45179_o;
  wire n45182_o;
  wire [7:0] n45187_o;
  wire n45190_o;
  wire [7:0] n45195_o;
  wire n45198_o;
  wire [7:0] n45203_o;
  wire n45206_o;
  wire [7:0] n45211_o;
  wire n45214_o;
  wire [7:0] n45219_o;
  wire n45226_o;
  wire n45228_o;
  wire n45230_o;
  wire n45232_o;
  wire n45234_o;
  wire n45236_o;
  wire n45238_o;
  wire n45240_o;
  wire n45242_o;
  wire [71:0] n45245_o;
  reg [5:0] n45246_q;
  wire [71:0] n45247_o;
  wire [7:0] n45248_data; // mem_rd
  wire [7:0] n45249_data; // mem_rd
  wire [7:0] n45250_data; // mem_rd
  wire [7:0] n45251_data; // mem_rd
  wire [7:0] n45252_data; // mem_rd
  wire [7:0] n45253_data; // mem_rd
  wire [7:0] n45254_data; // mem_rd
  wire [7:0] n45255_data; // mem_rd
  wire [7:0] n45256_data; // mem_rd
  wire [71:0] n45257_o;
  assign q_b = n45247_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:55:8  */
  assign q = n45257_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:56:8  */
  assign data = n45245_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:57:8  */
  assign address_r = n45246_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45129_o = q[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45130_o = q[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45131_o = q[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45132_o = q[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45133_o = q[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45134_o = q[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45135_o = q[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45136_o = q[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n45137_o = q[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45138_o = data_a[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45139_o = data_a[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45140_o = data_a[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45141_o = data_a[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45142_o = data_a[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45143_o = data_a[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45144_o = data_a[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45145_o = data_a[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n45146_o = data_a[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45150_o = byteena_a[0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45155_o = data[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45158_o = byteena_a[1];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45163_o = data[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45166_o = byteena_a[2];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45171_o = data[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45174_o = byteena_a[3];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45179_o = data[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45182_o = byteena_a[4];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45187_o = data[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45190_o = byteena_a[5];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45195_o = data[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45198_o = byteena_a[6];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45203_o = data[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45206_o = byteena_a[7];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45211_o = data[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n45214_o = byteena_a[8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n45219_o = data[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45226_o = wren_a & n45214_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45228_o = wren_a & n45206_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45230_o = wren_a & n45198_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45232_o = wren_a & n45190_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45234_o = wren_a & n45182_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45236_o = wren_a & n45174_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45238_o = wren_a & n45166_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45240_o = wren_a & n45158_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n45242_o = wren_a & n45150_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n45245_o = {n45138_o, n45139_o, n45140_o, n45141_o, n45142_o, n45143_o, n45144_o, n45145_o, n45146_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  always @(posedge clock0)
    n45246_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n45247_o = {n45137_o, n45136_o, n45135_o, n45134_o, n45133_o, n45132_o, n45131_o, n45130_o, n45129_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n1[63:0] ; // memory
  assign n45248_data = ram_block_n1[address_r];
  always @(posedge clock0)
    if (n45226_o)
      ram_block_n1[address_a] <= n45219_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n2[63:0] ; // memory
  assign n45249_data = ram_block_n2[address_r];
  always @(posedge clock0)
    if (n45228_o)
      ram_block_n2[address_a] <= n45211_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n3[63:0] ; // memory
  assign n45250_data = ram_block_n3[address_r];
  always @(posedge clock0)
    if (n45230_o)
      ram_block_n3[address_a] <= n45203_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n4[63:0] ; // memory
  assign n45251_data = ram_block_n4[address_r];
  always @(posedge clock0)
    if (n45232_o)
      ram_block_n4[address_a] <= n45195_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n5[63:0] ; // memory
  assign n45252_data = ram_block_n5[address_r];
  always @(posedge clock0)
    if (n45234_o)
      ram_block_n5[address_a] <= n45187_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n6[63:0] ; // memory
  assign n45253_data = ram_block_n6[address_r];
  always @(posedge clock0)
    if (n45236_o)
      ram_block_n6[address_a] <= n45179_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n7[63:0] ; // memory
  assign n45254_data = ram_block_n7[address_r];
  always @(posedge clock0)
    if (n45238_o)
      ram_block_n7[address_a] <= n45171_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n8[63:0] ; // memory
  assign n45255_data = ram_block_n8[address_r];
  always @(posedge clock0)
    if (n45240_o)
      ram_block_n8[address_a] <= n45163_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n9[63:0] ; // memory
  assign n45256_data = ram_block_n9[address_r];
  always @(posedge clock0)
    if (n45242_o)
      ram_block_n9[address_a] <= n45155_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  assign n45257_o = {n45256_data, n45255_data, n45254_data, n45253_data, n45252_data, n45251_data, n45250_data, n45249_data, n45248_data};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
endmodule

module sync_latch_72
  (input  enable_in,
   input  [71:0] data_in,
   output [71:0] data_out);
  wire [71:0] data_r;
  wire [71:0] n45121_o;
  assign data_out = data_r;
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:39:10  */
  assign data_r = n45121_o; // (signal)
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:45:4  */
  assign n45121_o = enable_in ? data_in : 72'b000000000000000000000000000000000000000000000000000000000000000000000000;
endmodule

module dpram_1024_1024_10_10_380_380
  (input  [9:0] address_a,
   input  clock,
   input  [379:0] data_a,
   input  wren_a,
   input  [9:0] address_b,
   output [379:0] q_b);
  wire [9:0] address_r;
  reg [9:0] n45114_q;
  wire [379:0] n45115_data; // mem_rd
  assign q_b = n45115_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n45114_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n45114_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [379:0] ram_block[1023:0] ; // memory
  assign n45115_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module ram2r1w_256_256_8_8_128_128
  (input  clock,
   input  clock_x2,
   input  [7:0] address_a,
   input  [15:0] byteena_a,
   input  [127:0] data_a,
   input  wren_a,
   input  [7:0] address1_b,
   input  [7:0] address2_b,
   output [127:0] q1_b,
   output [127:0] q2_b);
  wire wren;
  wire [7:0] address2_r;
  wire [7:0] address;
  wire [127:0] q_b;
  wire [127:0] q_latch;
  wire [7:0] address_a_r;
  wire [15:0] byteena_a_r;
  wire [127:0] data_a_r;
  reg wren_a_r;
  wire n45071_o;
  wire n45072_o;
  wire [7:0] n45073_o;
  wire [127:0] sync_latch_i_n45083;
  wire [127:0] sync_latch_i_data_out;
  wire [127:0] ram2_i_n45086;
  wire [127:0] ram2_i_q_b;
  reg [7:0] n45089_q;
  reg [7:0] n45090_q;
  reg [15:0] n45091_q;
  reg [127:0] n45092_q;
  reg n45093_q;
  assign q1_b = q_latch;
  assign q2_b = q_b;
  /* ../../HW/src/util/ram2r1w.vhd:71:8  */
  assign wren = n45071_o; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:72:8  */
  assign address2_r = n45089_q; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:73:8  */
  assign address = n45073_o; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:74:8  */
  assign q_b = ram2_i_n45086; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:75:8  */
  assign q_latch = sync_latch_i_n45083; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:76:8  */
  assign address_a_r = n45090_q; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:77:8  */
  assign byteena_a_r = n45091_q; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:78:8  */
  assign data_a_r = n45092_q; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:79:8  */
  always @*
    wren_a_r = n45093_q; // (isignal)
  initial
    wren_a_r = 1'b0;
  /* ../../HW/src/util/ram2r1w.vhd:85:18  */
  assign n45071_o = wren_a_r & clock;
  /* ../../HW/src/util/ram2r1w.vhd:86:33  */
  assign n45072_o = ~clock;
  /* ../../HW/src/util/ram2r1w.vhd:86:23  */
  assign n45073_o = n45072_o ? address1_b : address2_r;
  /* ../../HW/src/util/ram2r1w.vhd:108:17  */
  assign sync_latch_i_n45083 = sync_latch_i_data_out; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:99:1  */
  sync_latch_128 sync_latch_i (
    .enable_in(clock),
    .data_in(q_b),
    .data_out(sync_latch_i_data_out));
  /* ../../HW/src/util/ram2r1w.vhd:127:16  */
  assign ram2_i_n45086 = ram2_i_q_b; // (signal)
  /* ../../HW/src/util/ram2r1w.vhd:111:1  */
  dpram_be_256_256_8_8_128_128 ram2_i (
    .address_a(address_a_r),
    .byteena_a(byteena_a_r),
    .clock0(clock_x2),
    .data_a(data_a_r),
    .wren_a(wren),
    .address_b(address),
    .q_b(ram2_i_q_b));
  /* ../../HW/src/util/ram2r1w.vhd:90:4  */
  always @(posedge clock)
    n45089_q <= address2_b;
  /* ../../HW/src/util/ram2r1w.vhd:90:4  */
  always @(posedge clock)
    n45090_q <= address_a;
  /* ../../HW/src/util/ram2r1w.vhd:90:4  */
  always @(posedge clock)
    n45091_q <= byteena_a;
  /* ../../HW/src/util/ram2r1w.vhd:90:4  */
  always @(posedge clock)
    n45092_q <= data_a;
  /* ../../HW/src/util/ram2r1w.vhd:90:4  */
  always @(posedge clock)
    n45093_q <= wren_a;
  initial
    n45093_q = 1'b0;
endmodule

module shift_left_l_4_13
  (input  [12:0] data_in,
   input  [3:0] distance_in,
   output [12:0] data_out);
  wire [12:0] \input ;
  wire [12:0] \output ;
  wire [30:0] n45066_o;
  wire [12:0] n45067_o;
  assign data_out = \output ;
  /* ../../HW/platform/simulation/SLL.vhd:40:10  */
  assign \input  = data_in; // (signal)
  /* ../../HW/platform/simulation/SLL.vhd:41:10  */
  assign \output  = n45067_o; // (signal)
  /* ../../HW/platform/simulation/SLL.vhd:44:58  */
  assign n45066_o = {27'b0, distance_in};  //  uext
  /* ../../HW/platform/simulation/SLL.vhd:44:30  */
  assign n45067_o = \input  << n45066_o;
endmodule

module shift_right_l_4_13
  (input  [12:0] data_in,
   input  [3:0] distance_in,
   output [12:0] data_out);
  wire [12:0] \input ;
  wire [12:0] \output ;
  wire [30:0] n45063_o;
  wire [12:0] n45064_o;
  assign data_out = \output ;
  /* ../../HW/platform/simulation/SRL.vhd:40:10  */
  assign \input  = data_in; // (signal)
  /* ../../HW/platform/simulation/SRL.vhd:41:10  */
  assign \output  = n45064_o; // (signal)
  /* ../../HW/platform/simulation/SRL.vhd:44:59  */
  assign n45063_o = {27'b0, distance_in};  //  uext
  /* ../../HW/platform/simulation/SRL.vhd:44:30  */
  assign n45064_o = \input  >> n45063_o;
endmodule

module shift_left_a_4_13
  (input  [12:0] data_in,
   input  [3:0] distance_in,
   output [12:0] data_out);
  wire [12:0] \input ;
  wire [12:0] \output ;
  wire [30:0] n45060_o;
  wire [12:0] n45061_o;
  assign data_out = \output ;
  /* ../../HW/platform/simulation/SLA.vhd:40:10  */
  assign \input  = data_in; // (signal)
  /* ../../HW/platform/simulation/SLA.vhd:41:10  */
  assign \output  = n45061_o; // (signal)
  /* ../../HW/platform/simulation/SLA.vhd:45:58  */
  assign n45060_o = {27'b0, distance_in};  //  uext
  /* ../../HW/platform/simulation/SLA.vhd:45:30  */
  assign n45061_o = \input  << n45060_o;
endmodule

module shift_right_a_4_13
  (input  [12:0] data_in,
   input  [3:0] distance_in,
   output [12:0] data_out);
  wire [12:0] \input ;
  wire [12:0] \output ;
  wire [30:0] n45057_o;
  wire [12:0] n45058_o;
  assign data_out = \output ;
  /* ../../HW/platform/simulation/SRA.vhd:40:10  */
  assign \input  = data_in; // (signal)
  /* ../../HW/platform/simulation/SRA.vhd:41:10  */
  assign \output  = n45058_o; // (signal)
  /* ../../HW/platform/simulation/SRA.vhd:44:57  */
  assign n45057_o = {27'b0, distance_in};  //  uext
  /* ../../HW/platform/simulation/SRA.vhd:44:30  */
  assign n45058_o = $signed(\input ) >> n45057_o;
endmodule

module shift_left_a_2_32
  (input  [31:0] data_in,
   input  [1:0] distance_in,
   output [31:0] data_out);
  wire [31:0] \input ;
  wire [31:0] \output ;
  wire [30:0] n45054_o;
  wire [31:0] n45055_o;
  assign data_out = \output ;
  /* ../../HW/platform/simulation/SLA.vhd:40:10  */
  assign \input  = data_in; // (signal)
  /* ../../HW/platform/simulation/SLA.vhd:41:10  */
  assign \output  = n45055_o; // (signal)
  /* ../../HW/platform/simulation/SLA.vhd:45:58  */
  assign n45054_o = {29'b0, distance_in};  //  uext
  /* ../../HW/platform/simulation/SLA.vhd:45:30  */
  assign n45055_o = \input  << n45054_o;
endmodule

module shift_right_a_2_32
  (input  [31:0] data_in,
   input  [1:0] distance_in,
   output [31:0] data_out);
  wire [31:0] \input ;
  wire [31:0] \output ;
  wire [30:0] n45051_o;
  wire [31:0] n45052_o;
  assign data_out = \output ;
  /* ../../HW/platform/simulation/SRA.vhd:40:10  */
  assign \input  = data_in; // (signal)
  /* ../../HW/platform/simulation/SRA.vhd:41:10  */
  assign \output  = n45052_o; // (signal)
  /* ../../HW/platform/simulation/SRA.vhd:44:57  */
  assign n45051_o = {29'b0, distance_in};  //  uext
  /* ../../HW/platform/simulation/SRA.vhd:44:30  */
  assign n45052_o = $signed(\input ) >> n45051_o;
endmodule

module ramw_32_32_5_5_144_144
  (input  clock,
   input  clock_x2,
   input  [4:0] address_a,
   input  [17:0] byteena_a,
   input  [143:0] data_a,
   input  wren_a,
   input  [4:0] address_b,
   output [143:0] q_b);
  wire [71:0] data;
  wire [71:0] data_r;
  wire [8:0] byteena;
  wire [8:0] byteena_r;
  wire [5:0] waddress;
  wire [4:0] waddress_r;
  wire [5:0] raddress;
  wire [4:0] raddress_r;
  wire [71:0] q;
  wire [71:0] q_latch;
  wire wren;
  wire wren_r;
  wire [71:0] n45009_o;
  wire n45010_o;
  wire [71:0] n45011_o;
  wire [8:0] n45012_o;
  wire n45013_o;
  wire [8:0] n45014_o;
  wire n45015_o;
  wire [4:0] n45016_o;
  wire n45017_o;
  wire n45018_o;
  wire [4:0] n45019_o;
  wire n45020_o;
  wire n45021_o;
  wire n45022_o;
  wire n45023_o;
  wire n45024_o;
  wire [71:0] sync_latch_i_n45025;
  wire [71:0] sync_latch_i_data_out;
  wire [71:0] n45031_o;
  wire [8:0] n45032_o;
  wire [71:0] ram_i_n45039;
  wire [71:0] ram_i_q_b;
  reg [71:0] n45042_q;
  reg [8:0] n45043_q;
  wire [5:0] n45044_o;
  reg [4:0] n45045_q;
  wire [5:0] n45046_o;
  reg [4:0] n45047_q;
  reg n45048_q;
  wire [143:0] n45049_o;
  assign q_b = n45049_o;
  /* ../../HW/src/util/ramw.vhd:55:8  */
  assign data = n45011_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:56:8  */
  assign data_r = n45042_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:57:8  */
  assign byteena = n45014_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:58:8  */
  assign byteena_r = n45043_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:59:8  */
  assign waddress = n45044_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:60:8  */
  assign waddress_r = n45045_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:61:8  */
  assign raddress = n45046_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:62:8  */
  assign raddress_r = n45047_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:63:8  */
  assign q = ram_i_n45039; // (signal)
  /* ../../HW/src/util/ramw.vhd:64:8  */
  assign q_latch = sync_latch_i_n45025; // (signal)
  /* ../../HW/src/util/ramw.vhd:65:8  */
  assign wren = n45024_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:66:8  */
  assign wren_r = n45048_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:69:15  */
  assign n45009_o = data_a[143:72];
  /* ../../HW/src/util/ramw.vhd:69:66  */
  assign n45010_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:69:56  */
  assign n45011_o = n45010_o ? n45009_o : data_r;
  /* ../../HW/src/util/ramw.vhd:70:21  */
  assign n45012_o = byteena_a[17:9];
  /* ../../HW/src/util/ramw.vhd:70:78  */
  assign n45013_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:70:68  */
  assign n45014_o = n45013_o ? n45012_o : byteena_r;
  /* ../../HW/src/util/ramw.vhd:71:61  */
  assign n45015_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:71:51  */
  assign n45016_o = n45015_o ? address_a : waddress_r;
  /* ../../HW/src/util/ramw.vhd:72:17  */
  assign n45017_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:73:61  */
  assign n45018_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:73:51  */
  assign n45019_o = n45018_o ? address_b : raddress_r;
  /* ../../HW/src/util/ramw.vhd:74:17  */
  assign n45020_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:77:17  */
  assign n45021_o = wren_r & clock;
  /* ../../HW/src/util/ramw.vhd:77:44  */
  assign n45022_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:77:39  */
  assign n45023_o = wren_a & n45022_o;
  /* ../../HW/src/util/ramw.vhd:77:28  */
  assign n45024_o = n45021_o | n45023_o;
  /* ../../HW/src/util/ramw.vhd:88:17  */
  assign sync_latch_i_n45025 = sync_latch_i_data_out; // (signal)
  /* ../../HW/src/util/ramw.vhd:79:1  */
  sync_latch_72 sync_latch_i (
    .enable_in(clock),
    .data_in(q),
    .data_out(sync_latch_i_data_out));
  /* ../../HW/src/util/ramw.vhd:94:23  */
  assign n45031_o = data_a[71:0];
  /* ../../HW/src/util/ramw.vhd:95:29  */
  assign n45032_o = byteena_a[8:0];
  /* ../../HW/src/util/ramw.vhd:116:14  */
  assign ram_i_n45039 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/ramw.vhd:102:1  */
  dpram_be_64_64_6_6_72_72 ram_i (
    .address_a(waddress),
    .byteena_a(byteena),
    .clock0(clock_x2),
    .data_a(data),
    .wren_a(wren),
    .address_b(raddress),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n45042_q <= n45031_o;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n45043_q <= n45032_o;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  assign n45044_o = {n45016_o, n45017_o};
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n45045_q <= address_a;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  assign n45046_o = {n45019_o, n45020_o};
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n45047_q <= address_b;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n45048_q <= wren_a;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  assign n45049_o = {q_latch, q};
endmodule

module dpram_be_512_512_9_9_136_136
  (input  [8:0] address_a,
   input  [16:0] byteena_a,
   input  clock0,
   input  [135:0] data_a,
   input  wren_a,
   input  [8:0] address_b,
   output [135:0] q_b);
  wire [135:0] q;
  wire [135:0] data;
  wire [8:0] address_r;
  wire [7:0] n44758_o;
  wire [7:0] n44759_o;
  wire [7:0] n44760_o;
  wire [7:0] n44761_o;
  wire [7:0] n44762_o;
  wire [7:0] n44763_o;
  wire [7:0] n44764_o;
  wire [7:0] n44765_o;
  wire [7:0] n44766_o;
  wire [7:0] n44767_o;
  wire [7:0] n44768_o;
  wire [7:0] n44769_o;
  wire [7:0] n44770_o;
  wire [7:0] n44771_o;
  wire [7:0] n44772_o;
  wire [7:0] n44773_o;
  wire [7:0] n44774_o;
  wire [7:0] n44775_o;
  wire [7:0] n44776_o;
  wire [7:0] n44777_o;
  wire [7:0] n44778_o;
  wire [7:0] n44779_o;
  wire [7:0] n44780_o;
  wire [7:0] n44781_o;
  wire [7:0] n44782_o;
  wire [7:0] n44783_o;
  wire [7:0] n44784_o;
  wire [7:0] n44785_o;
  wire [7:0] n44786_o;
  wire [7:0] n44787_o;
  wire [7:0] n44788_o;
  wire [7:0] n44789_o;
  wire [7:0] n44790_o;
  wire [7:0] n44791_o;
  wire n44795_o;
  wire [7:0] n44800_o;
  wire n44803_o;
  wire [7:0] n44808_o;
  wire n44811_o;
  wire [7:0] n44816_o;
  wire n44819_o;
  wire [7:0] n44824_o;
  wire n44827_o;
  wire [7:0] n44832_o;
  wire n44835_o;
  wire [7:0] n44840_o;
  wire n44843_o;
  wire [7:0] n44848_o;
  wire n44851_o;
  wire [7:0] n44856_o;
  wire n44859_o;
  wire [7:0] n44864_o;
  wire n44867_o;
  wire [7:0] n44872_o;
  wire n44875_o;
  wire [7:0] n44880_o;
  wire n44883_o;
  wire [7:0] n44888_o;
  wire n44891_o;
  wire [7:0] n44896_o;
  wire n44899_o;
  wire [7:0] n44904_o;
  wire n44907_o;
  wire [7:0] n44912_o;
  wire n44915_o;
  wire [7:0] n44920_o;
  wire n44923_o;
  wire [7:0] n44928_o;
  wire n44935_o;
  wire n44937_o;
  wire n44939_o;
  wire n44941_o;
  wire n44943_o;
  wire n44945_o;
  wire n44947_o;
  wire n44949_o;
  wire n44951_o;
  wire n44953_o;
  wire n44955_o;
  wire n44957_o;
  wire n44959_o;
  wire n44961_o;
  wire n44963_o;
  wire n44965_o;
  wire n44967_o;
  wire [135:0] n44970_o;
  reg [8:0] n44971_q;
  wire [135:0] n44972_o;
  wire [7:0] n44973_data; // mem_rd
  wire [7:0] n44974_data; // mem_rd
  wire [7:0] n44975_data; // mem_rd
  wire [7:0] n44976_data; // mem_rd
  wire [7:0] n44977_data; // mem_rd
  wire [7:0] n44978_data; // mem_rd
  wire [7:0] n44979_data; // mem_rd
  wire [7:0] n44980_data; // mem_rd
  wire [7:0] n44981_data; // mem_rd
  wire [7:0] n44982_data; // mem_rd
  wire [7:0] n44983_data; // mem_rd
  wire [7:0] n44984_data; // mem_rd
  wire [7:0] n44985_data; // mem_rd
  wire [7:0] n44986_data; // mem_rd
  wire [7:0] n44987_data; // mem_rd
  wire [7:0] n44988_data; // mem_rd
  wire [7:0] n44989_data; // mem_rd
  wire [135:0] n44990_o;
  assign q_b = n44972_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:55:8  */
  assign q = n44990_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:56:8  */
  assign data = n44970_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:57:8  */
  assign address_r = n44971_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44758_o = q[135:128];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44759_o = q[127:120];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44760_o = q[119:112];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44761_o = q[111:104];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44762_o = q[103:96];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44763_o = q[95:88];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44764_o = q[87:80];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44765_o = q[79:72];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44766_o = q[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44767_o = q[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44768_o = q[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44769_o = q[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44770_o = q[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44771_o = q[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44772_o = q[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44773_o = q[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n44774_o = q[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44775_o = data_a[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44776_o = data_a[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44777_o = data_a[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44778_o = data_a[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44779_o = data_a[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44780_o = data_a[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44781_o = data_a[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44782_o = data_a[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44783_o = data_a[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44784_o = data_a[79:72];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44785_o = data_a[87:80];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44786_o = data_a[95:88];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44787_o = data_a[103:96];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44788_o = data_a[111:104];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44789_o = data_a[119:112];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44790_o = data_a[127:120];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n44791_o = data_a[135:128];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44795_o = byteena_a[0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44800_o = data[135:128];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44803_o = byteena_a[1];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44808_o = data[127:120];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44811_o = byteena_a[2];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44816_o = data[119:112];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44819_o = byteena_a[3];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44824_o = data[111:104];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44827_o = byteena_a[4];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44832_o = data[103:96];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44835_o = byteena_a[5];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44840_o = data[95:88];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44843_o = byteena_a[6];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44848_o = data[87:80];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44851_o = byteena_a[7];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44856_o = data[79:72];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44859_o = byteena_a[8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44864_o = data[71:64];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44867_o = byteena_a[9];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44872_o = data[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44875_o = byteena_a[10];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44880_o = data[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44883_o = byteena_a[11];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44888_o = data[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44891_o = byteena_a[12];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44896_o = data[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44899_o = byteena_a[13];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44904_o = data[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44907_o = byteena_a[14];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44912_o = data[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44915_o = byteena_a[15];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44920_o = data[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n44923_o = byteena_a[16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n44928_o = data[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44935_o = wren_a & n44923_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44937_o = wren_a & n44915_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44939_o = wren_a & n44907_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44941_o = wren_a & n44899_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44943_o = wren_a & n44891_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44945_o = wren_a & n44883_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44947_o = wren_a & n44875_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44949_o = wren_a & n44867_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44951_o = wren_a & n44859_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44953_o = wren_a & n44851_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44955_o = wren_a & n44843_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44957_o = wren_a & n44835_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44959_o = wren_a & n44827_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44961_o = wren_a & n44819_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44963_o = wren_a & n44811_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44965_o = wren_a & n44803_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n44967_o = wren_a & n44795_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n44970_o = {n44775_o, n44776_o, n44777_o, n44778_o, n44779_o, n44780_o, n44781_o, n44782_o, n44783_o, n44784_o, n44785_o, n44786_o, n44787_o, n44788_o, n44789_o, n44790_o, n44791_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  always @(posedge clock0)
    n44971_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n44972_o = {n44774_o, n44773_o, n44772_o, n44771_o, n44770_o, n44769_o, n44768_o, n44767_o, n44766_o, n44765_o, n44764_o, n44763_o, n44762_o, n44761_o, n44760_o, n44759_o, n44758_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n1[511:0] ; // memory
  assign n44973_data = ram_block_n1[address_r];
  always @(posedge clock0)
    if (n44935_o)
      ram_block_n1[address_a] <= n44928_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n2[511:0] ; // memory
  assign n44974_data = ram_block_n2[address_r];
  always @(posedge clock0)
    if (n44937_o)
      ram_block_n2[address_a] <= n44920_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n3[511:0] ; // memory
  assign n44975_data = ram_block_n3[address_r];
  always @(posedge clock0)
    if (n44939_o)
      ram_block_n3[address_a] <= n44912_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n4[511:0] ; // memory
  assign n44976_data = ram_block_n4[address_r];
  always @(posedge clock0)
    if (n44941_o)
      ram_block_n4[address_a] <= n44904_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n5[511:0] ; // memory
  assign n44977_data = ram_block_n5[address_r];
  always @(posedge clock0)
    if (n44943_o)
      ram_block_n5[address_a] <= n44896_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n6[511:0] ; // memory
  assign n44978_data = ram_block_n6[address_r];
  always @(posedge clock0)
    if (n44945_o)
      ram_block_n6[address_a] <= n44888_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n7[511:0] ; // memory
  assign n44979_data = ram_block_n7[address_r];
  always @(posedge clock0)
    if (n44947_o)
      ram_block_n7[address_a] <= n44880_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n8[511:0] ; // memory
  assign n44980_data = ram_block_n8[address_r];
  always @(posedge clock0)
    if (n44949_o)
      ram_block_n8[address_a] <= n44872_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n9[511:0] ; // memory
  assign n44981_data = ram_block_n9[address_r];
  always @(posedge clock0)
    if (n44951_o)
      ram_block_n9[address_a] <= n44864_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n10[511:0] ; // memory
  assign n44982_data = ram_block_n10[address_r];
  always @(posedge clock0)
    if (n44953_o)
      ram_block_n10[address_a] <= n44856_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n11[511:0] ; // memory
  assign n44983_data = ram_block_n11[address_r];
  always @(posedge clock0)
    if (n44955_o)
      ram_block_n11[address_a] <= n44848_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n12[511:0] ; // memory
  assign n44984_data = ram_block_n12[address_r];
  always @(posedge clock0)
    if (n44957_o)
      ram_block_n12[address_a] <= n44840_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n13[511:0] ; // memory
  assign n44985_data = ram_block_n13[address_r];
  always @(posedge clock0)
    if (n44959_o)
      ram_block_n13[address_a] <= n44832_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n14[511:0] ; // memory
  assign n44986_data = ram_block_n14[address_r];
  always @(posedge clock0)
    if (n44961_o)
      ram_block_n14[address_a] <= n44824_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n15[511:0] ; // memory
  assign n44987_data = ram_block_n15[address_r];
  always @(posedge clock0)
    if (n44963_o)
      ram_block_n15[address_a] <= n44816_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n16[511:0] ; // memory
  assign n44988_data = ram_block_n16[address_r];
  always @(posedge clock0)
    if (n44965_o)
      ram_block_n16[address_a] <= n44808_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n17[511:0] ; // memory
  assign n44989_data = ram_block_n17[address_r];
  always @(posedge clock0)
    if (n44967_o)
      ram_block_n17[address_a] <= n44800_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  assign n44990_o = {n44989_data, n44988_data, n44987_data, n44986_data, n44985_data, n44984_data, n44983_data, n44982_data, n44981_data, n44980_data, n44979_data, n44978_data, n44977_data, n44976_data, n44975_data, n44974_data, n44973_data};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
endmodule

module sync_latch_136
  (input  enable_in,
   input  [135:0] data_in,
   output [135:0] data_out);
  wire [135:0] data_r;
  wire [135:0] n44750_o;
  assign data_out = data_r;
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:39:10  */
  assign data_r = n44750_o; // (signal)
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:45:4  */
  assign n44750_o = enable_in ? data_in : 136'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endmodule

module scfifo_380_10_4_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [379:0] data_in,
   input  write_in,
   input  read_in,
   output [379:0] q_out,
   output [9:0] ravail_out,
   output [9:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [379:0] q;
  wire [9:0] address_a;
  wire [9:0] address_b;
  wire [9:0] waddr_r;
  wire [9:0] waddr_rr;
  wire [9:0] raddr_r;
  wire [9:0] raddr;
  wire [9:0] ravail;
  wire [9:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [379:0] ram_i_n44679;
  wire [379:0] ram_i_q_b;
  wire [9:0] n44682_o;
  wire [9:0] n44683_o;
  wire n44684_o;
  wire n44687_o;
  wire n44688_o;
  wire [9:0] n44691_o;
  wire [9:0] n44692_o;
  wire n44695_o;
  wire [9:0] n44698_o;
  wire [9:0] n44700_o;
  wire n44701_o;
  wire n44704_o;
  wire [9:0] n44706_o;
  wire n44707_o;
  wire n44710_o;
  wire n44712_o;
  wire n44714_o;
  wire n44717_o;
  wire [9:0] n44739_o;
  reg [9:0] n44740_q;
  reg [9:0] n44741_q;
  reg [9:0] n44742_q;
  reg n44744_q;
  reg n44745_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n44684_o;
  assign full_out = full_r;
  assign almost_full_out = n44688_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n44679; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n44740_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n44741_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n44742_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n44692_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n44682_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n44683_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n44744_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n44745_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n44679 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_1024_1024_10_10_380_380 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n44682_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n44683_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n44684_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n44687_o = $unsigned(wused) >= $unsigned(10'b0000000100);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n44688_o = n44687_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n44691_o = raddr_r + 10'b0000000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n44692_o = read_in ? n44691_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n44695_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n44698_o = waddr_r + 10'b0000000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n44700_o = waddr_r + 10'b0000000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n44701_o = n44700_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n44704_o = n44701_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n44706_o = waddr_r + 10'b0000000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n44707_o = n44706_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n44710_o = n44707_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n44712_o = write_in ? n44704_o : n44710_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n44714_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n44717_o = n44714_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n44739_o = write_in ? n44698_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n44695_o)
    if (n44695_o)
      n44740_q <= 10'b0000000000;
    else
      n44740_q <= n44739_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n44695_o)
    if (n44695_o)
      n44741_q <= 10'b0000000000;
    else
      n44741_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n44695_o)
    if (n44695_o)
      n44742_q <= 10'b0000000000;
    else
      n44742_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n44695_o)
    if (n44695_o)
      n44744_q <= 1'b0;
    else
      n44744_q <= n44717_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n44695_o)
    if (n44695_o)
      n44745_q <= 1'b0;
    else
      n44745_q <= n44712_o;
endmodule

module delayv_8_6
  (input  clock_in,
   input  reset_in,
   input  [7:0] in_in,
   input  enable_in,
   output [7:0] out_out);
  wire [47:0] fifo_r;
  wire [7:0] n44639_o;
  wire n44642_o;
  wire [7:0] n44650_o;
  wire [7:0] n44651_o;
  wire [7:0] n44652_o;
  wire [7:0] n44653_o;
  wire [7:0] n44654_o;
  wire [7:0] n44655_o;
  wire [7:0] n44656_o;
  wire [7:0] n44657_o;
  wire [7:0] n44658_o;
  wire [7:0] n44659_o;
  wire [7:0] n44660_o;
  wire [7:0] n44661_o;
  wire [7:0] n44662_o;
  wire [7:0] n44663_o;
  wire [7:0] n44664_o;
  wire [7:0] n44665_o;
  wire [7:0] n44666_o;
  wire [47:0] n44667_o;
  wire [47:0] n44669_o;
  reg [47:0] n44672_q;
  assign out_out = n44639_o;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n44672_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:48:18  */
  assign n44639_o = fifo_r[7:0];
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n44642_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44650_o = fifo_r[15:8];
  assign n44651_o = fifo_r[7:0];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44652_o = enable_in ? n44650_o : n44651_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44653_o = fifo_r[23:16];
  assign n44654_o = fifo_r[15:8];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44655_o = enable_in ? n44653_o : n44654_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44656_o = fifo_r[31:24];
  assign n44657_o = fifo_r[23:16];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44658_o = enable_in ? n44656_o : n44657_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44659_o = fifo_r[39:32];
  assign n44660_o = fifo_r[31:24];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44661_o = enable_in ? n44659_o : n44660_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44662_o = fifo_r[47:40];
  assign n44663_o = fifo_r[39:32];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44664_o = enable_in ? n44662_o : n44663_o;
  assign n44665_o = fifo_r[47:40];
  /* ../../HW/src/util/delayv.vhd:64:13  */
  assign n44666_o = enable_in ? in_in : n44665_o;
  assign n44667_o = {n44666_o, n44664_o, n44661_o, n44658_o, n44655_o, n44652_o};
  assign n44669_o = {8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000, 8'b00000000};
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n44642_o)
    if (n44642_o)
      n44672_q <= n44669_o;
    else
      n44672_q <= n44667_o;
endmodule

module delayv_12_6
  (input  clock_in,
   input  reset_in,
   input  [11:0] in_in,
   input  enable_in,
   output [11:0] out_out);
  wire [71:0] fifo_r;
  wire [11:0] n44604_o;
  wire n44607_o;
  wire [11:0] n44615_o;
  wire [11:0] n44616_o;
  wire [11:0] n44617_o;
  wire [11:0] n44618_o;
  wire [11:0] n44619_o;
  wire [11:0] n44620_o;
  wire [11:0] n44621_o;
  wire [11:0] n44622_o;
  wire [11:0] n44623_o;
  wire [11:0] n44624_o;
  wire [11:0] n44625_o;
  wire [11:0] n44626_o;
  wire [11:0] n44627_o;
  wire [11:0] n44628_o;
  wire [11:0] n44629_o;
  wire [11:0] n44630_o;
  wire [11:0] n44631_o;
  wire [71:0] n44632_o;
  wire [71:0] n44634_o;
  reg [71:0] n44637_q;
  assign out_out = n44604_o;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n44637_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:48:18  */
  assign n44604_o = fifo_r[11:0];
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n44607_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44615_o = fifo_r[23:12];
  assign n44616_o = fifo_r[11:0];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44617_o = enable_in ? n44615_o : n44616_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44618_o = fifo_r[35:24];
  assign n44619_o = fifo_r[23:12];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44620_o = enable_in ? n44618_o : n44619_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44621_o = fifo_r[47:36];
  assign n44622_o = fifo_r[35:24];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44623_o = enable_in ? n44621_o : n44622_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44624_o = fifo_r[59:48];
  assign n44625_o = fifo_r[47:36];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44626_o = enable_in ? n44624_o : n44625_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n44627_o = fifo_r[71:60];
  assign n44628_o = fifo_r[59:48];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n44629_o = enable_in ? n44627_o : n44628_o;
  assign n44630_o = fifo_r[71:60];
  /* ../../HW/src/util/delayv.vhd:64:13  */
  assign n44631_o = enable_in ? in_in : n44630_o;
  assign n44632_o = {n44631_o, n44629_o, n44626_o, n44623_o, n44620_o, n44617_o};
  assign n44634_o = {12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000};
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n44607_o)
    if (n44607_o)
      n44637_q <= n44634_o;
    else
      n44637_q <= n44632_o;
endmodule

module delayv_8_1
  (input  clock_in,
   input  reset_in,
   input  [7:0] in_in,
   input  enable_in,
   output [7:0] out_out);
  wire [7:0] fifo_r;
  wire n44594_o;
  wire [7:0] n44601_o;
  reg [7:0] n44602_q;
  assign out_out = fifo_r;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n44602_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n44594_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:56:9  */
  assign n44601_o = enable_in ? in_in : fifo_r;
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n44594_o)
    if (n44594_o)
      n44602_q <= 8'b00000000;
    else
      n44602_q <= n44601_o;
endmodule

module delay_6
  (input  clock_in,
   input  reset_in,
   input  in_in,
   input  enable_in,
   output out_out);
  wire [5:0] fifo_r;
  wire n44557_o;
  wire n44560_o;
  wire n44568_o;
  wire n44569_o;
  wire n44570_o;
  wire n44571_o;
  wire n44572_o;
  wire n44573_o;
  wire n44574_o;
  wire n44575_o;
  wire n44576_o;
  wire n44577_o;
  wire n44578_o;
  wire n44579_o;
  wire n44580_o;
  wire n44581_o;
  wire n44582_o;
  wire n44583_o;
  wire n44584_o;
  wire [5:0] n44585_o;
  wire [5:0] n44587_o;
  reg [5:0] n44590_q;
  assign out_out = n44557_o;
  /* ../../HW/src/util/delay.vhd:46:8  */
  assign fifo_r = n44590_q; // (signal)
  /* ../../HW/src/util/delay.vhd:48:18  */
  assign n44557_o = fifo_r[0];
  /* ../../HW/src/util/delay.vhd:51:16  */
  assign n44560_o = ~reset_in;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n44568_o = fifo_r[1];
  /* ../../HW/src/pcore/register_file.vhd:231:1  */
  assign n44569_o = fifo_r[0];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n44570_o = enable_in ? n44568_o : n44569_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n44571_o = fifo_r[2];
  assign n44572_o = fifo_r[1];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n44573_o = enable_in ? n44571_o : n44572_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n44574_o = fifo_r[3];
  /* ../../HW/src/pcore/register_file.vhd:193:10  */
  assign n44575_o = fifo_r[2];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n44576_o = enable_in ? n44574_o : n44575_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n44577_o = fifo_r[4];
  /* ../../HW/src/pcore/register_file.vhd:233:4  */
  assign n44578_o = fifo_r[3];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n44579_o = enable_in ? n44577_o : n44578_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n44580_o = fifo_r[5];
  assign n44581_o = fifo_r[4];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n44582_o = enable_in ? n44580_o : n44581_o;
  assign n44583_o = fifo_r[5];
  /* ../../HW/src/util/delay.vhd:64:13  */
  assign n44584_o = enable_in ? in_in : n44583_o;
  assign n44585_o = {n44584_o, n44582_o, n44579_o, n44576_o, n44573_o, n44570_o};
  assign n44587_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/util/delay.vhd:56:9  */
  always @(posedge clock_in or posedge n44560_o)
    if (n44560_o)
      n44590_q <= n44587_o;
    else
      n44590_q <= n44585_o;
endmodule

module register_file
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  rd_en_in,
   input  rd_x1_vector_in,
   input  [11:0] rd_x1_addr_in,
   input  rd_x2_vector_in,
   input  [11:0] rd_x2_addr_in,
   input  wr_en_in,
   input  wr_vector_in,
   input  [11:0] wr_addr_in,
   input  [95:0] wr_data_in,
   input  [7:0] wr_lane_in,
   input  [2:0] dp_rd_vector_in,
   input  [1:0] dp_rd_scatter_in,
   input  [2:0] dp_rd_scatter_cnt_in,
   input  [2:0] dp_rd_scatter_vector_in,
   input  dp_rd_gen_valid_in,
   input  [1:0] dp_rd_data_flow_in,
   input  [1:0] dp_rd_data_type_in,
   input  dp_rd_stream_in,
   input  [1:0] dp_rd_stream_id_in,
   input  [16:0] dp_rd_addr_in,
   input  [2:0] dp_wr_vector_in,
   input  [16:0] dp_wr_addr_in,
   input  dp_write_in,
   input  dp_read_in,
   input  [95:0] dp_writedata_in,
   output rd_en_out,
   output [95:0] rd_x1_data_out,
   output [95:0] rd_x2_data_out,
   output [95:0] dp_readdata_out,
   output dp_readena_out);
  wire [7:0] wr_lane;
  wire [8:0] rd_x1_addr;
  wire [8:0] rd_x2_addr;
  wire [8:0] wr_addr;
  wire [95:0] wr_data;
  wire [95:0] wr_data2;
  wire wr_en;
  wire rd_en_r;
  wire rd_en_rr;
  wire [95:0] q1;
  wire [95:0] q2;
  wire dp_rd_en_r;
  wire dp_rd_en_rr;
  wire [2:0] wr_vaddr;
  wire [2:0] wr_vector;
  wire [15:0] byteena;
  wire [16:0] dp_rd_addr;
  wire [16:0] dp_wr_addr;
  wire [95:0] dp_writedata;
  wire [127:0] wr_data2_ram;
  wire [127:0] q1_ram;
  wire [127:0] q1_ram_r;
  wire [127:0] q2_ram;
  wire [127:0] q2_ram_r;
  wire n44342_o;
  wire n44343_o;
  wire [8:0] n44345_o;
  wire [8:0] n44346_o;
  wire [8:0] n44347_o;
  wire [2:0] n44348_o;
  wire [2:0] n44349_o;
  wire [2:0] n44350_o;
  wire [95:0] n44351_o;
  wire [2:0] n44352_o;
  wire [2:0] n44353_o;
  wire [7:0] n44354_o;
  wire [8:0] n44356_o;
  wire [8:0] n44357_o;
  wire [8:0] n44358_o;
  wire [8:0] n44359_o;
  wire n44364_o;
  wire n44365_o;
  wire n44366_o;
  wire [1:0] n44367_o;
  wire n44368_o;
  wire n44369_o;
  wire [1:0] n44370_o;
  wire n44371_o;
  wire n44372_o;
  wire [1:0] n44373_o;
  wire n44374_o;
  wire n44375_o;
  wire [1:0] n44376_o;
  wire n44377_o;
  wire n44378_o;
  wire [1:0] n44379_o;
  wire n44380_o;
  wire n44381_o;
  wire [1:0] n44382_o;
  wire n44383_o;
  wire n44384_o;
  wire [1:0] n44385_o;
  wire n44386_o;
  wire n44387_o;
  wire [1:0] n44388_o;
  wire [2:0] n44389_o;
  wire [2:0] n44391_o;
  wire [2:0] n44392_o;
  wire n44393_o;
  wire [1:0] n44396_o;
  wire [2:0] n44398_o;
  wire [2:0] n44399_o;
  wire n44400_o;
  wire [1:0] n44403_o;
  wire [2:0] n44405_o;
  wire [2:0] n44406_o;
  wire n44407_o;
  wire [1:0] n44410_o;
  wire [2:0] n44412_o;
  wire [2:0] n44413_o;
  wire n44414_o;
  wire [1:0] n44417_o;
  wire [2:0] n44419_o;
  wire [2:0] n44420_o;
  wire n44421_o;
  wire [1:0] n44424_o;
  wire [2:0] n44426_o;
  wire [2:0] n44427_o;
  wire n44428_o;
  wire [1:0] n44431_o;
  wire [2:0] n44433_o;
  wire [2:0] n44434_o;
  wire n44435_o;
  wire [1:0] n44438_o;
  wire [2:0] n44440_o;
  wire [2:0] n44441_o;
  wire n44442_o;
  wire [1:0] n44445_o;
  wire [15:0] n44446_o;
  wire [15:0] n44447_o;
  wire [15:0] n44448_o;
  wire n44454_o;
  wire [11:0] n44455_o;
  wire [11:0] n44456_o;
  wire [23:0] n44457_o;
  wire [11:0] n44458_o;
  wire [35:0] n44459_o;
  wire [11:0] n44460_o;
  wire [47:0] n44461_o;
  wire [11:0] n44462_o;
  wire [59:0] n44463_o;
  wire [11:0] n44464_o;
  wire [71:0] n44465_o;
  wire [11:0] n44466_o;
  wire [83:0] n44467_o;
  wire [11:0] n44468_o;
  wire [95:0] n44469_o;
  wire [95:0] n44470_o;
  wire n44474_o;
  wire [11:0] n44492_o;
  wire [11:0] n44493_o;
  wire [11:0] n44494_o;
  wire [11:0] n44496_o;
  wire [11:0] n44497_o;
  wire [11:0] n44498_o;
  wire [11:0] n44500_o;
  wire [11:0] n44501_o;
  wire [11:0] n44502_o;
  wire [11:0] n44504_o;
  wire [11:0] n44505_o;
  wire [11:0] n44506_o;
  wire [11:0] n44508_o;
  wire [11:0] n44509_o;
  wire [11:0] n44510_o;
  wire [11:0] n44512_o;
  wire [11:0] n44513_o;
  wire [11:0] n44514_o;
  wire [11:0] n44516_o;
  wire [11:0] n44517_o;
  wire [11:0] n44518_o;
  wire [11:0] n44520_o;
  wire [11:0] n44521_o;
  wire [11:0] n44522_o;
  wire n44526_o;
  wire n44530_o;
  wire [7:0] n44538_o;
  wire [7:0] n44539_o;
  wire [127:0] ram3_i_n44540;
  wire [7:0] n44541_o;
  wire [127:0] ram3_i_n44542;
  wire [127:0] ram3_i_q1_b;
  wire [127:0] ram3_i_q2_b;
  reg n44547_q;
  reg n44548_q;
  wire [95:0] n44549_o;
  wire [95:0] n44550_o;
  reg n44551_q;
  reg n44552_q;
  wire [127:0] n44553_o;
  reg [127:0] n44554_q;
  reg [127:0] n44555_q;
  assign rd_en_out = rd_en_rr;
  assign rd_x1_data_out = q1;
  assign rd_x2_data_out = q2;
  assign dp_readdata_out = q2;
  assign dp_readena_out = dp_rd_en_rr;
  /* ../../HW/src/pcore/register_file.vhd:84:8  */
  assign wr_lane = n44354_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:85:8  */
  assign rd_x1_addr = n44356_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:86:8  */
  assign rd_x2_addr = n44358_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:87:8  */
  assign wr_addr = n44346_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:88:8  */
  assign wr_data = n44351_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:89:8  */
  assign wr_data2 = n44470_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:90:8  */
  assign wr_en = n44343_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:91:8  */
  assign rd_en_r = n44547_q; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:92:8  */
  assign rd_en_rr = n44548_q; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:93:8  */
  assign q1 = n44549_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:94:8  */
  assign q2 = n44550_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:95:8  */
  assign dp_rd_en_r = n44551_q; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:96:8  */
  assign dp_rd_en_rr = n44552_q; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:97:8  */
  assign wr_vaddr = n44349_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:99:8  */
  assign wr_vector = n44353_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:100:8  */
  assign byteena = n44448_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:102:8  */
  assign dp_rd_addr = dp_rd_addr_in; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:103:8  */
  assign dp_wr_addr = dp_wr_addr_in; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:105:8  */
  assign dp_writedata = dp_writedata_in; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:107:8  */
  assign wr_data2_ram = n44553_o; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:108:8  */
  assign q1_ram = ram3_i_n44540; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:109:8  */
  assign q1_ram_r = n44554_q; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:110:8  */
  assign q2_ram = ram3_i_n44542; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:111:8  */
  assign q2_ram_r = n44555_q; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:166:36  */
  assign n44342_o = dp_write_in | wr_en_in;
  /* ../../HW/src/pcore/register_file.vhd:166:14  */
  assign n44343_o = n44342_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/register_file.vhd:168:22  */
  assign n44345_o = wr_addr_in[11:3];
  /* ../../HW/src/pcore/register_file.vhd:168:70  */
  assign n44346_o = wr_en_in ? n44345_o : n44347_o;
  /* ../../HW/src/pcore/register_file.vhd:168:105  */
  assign n44347_o = dp_wr_addr[11:3];
  /* ../../HW/src/pcore/register_file.vhd:170:23  */
  assign n44348_o = wr_addr_in[2:0];
  /* ../../HW/src/pcore/register_file.vhd:170:51  */
  assign n44349_o = wr_en_in ? n44348_o : n44350_o;
  /* ../../HW/src/pcore/register_file.vhd:170:86  */
  assign n44350_o = dp_wr_addr[2:0];
  /* ../../HW/src/pcore/register_file.vhd:172:23  */
  assign n44351_o = wr_en_in ? wr_data_in : dp_writedata;
  assign n44352_o = {wr_vector_in, wr_vector_in, wr_vector_in};
  /* ../../HW/src/pcore/register_file.vhd:174:37  */
  assign n44353_o = wr_en_in ? n44352_o : dp_wr_vector_in;
  /* ../../HW/src/pcore/register_file.vhd:176:23  */
  assign n44354_o = wr_en_in ? wr_lane_in : 8'b11111111;
  /* ../../HW/src/pcore/register_file.vhd:180:28  */
  assign n44356_o = rd_x1_addr_in[11:3];
  /* ../../HW/src/pcore/register_file.vhd:182:28  */
  assign n44357_o = rd_x2_addr_in[11:3];
  /* ../../HW/src/pcore/register_file.vhd:182:76  */
  assign n44358_o = rd_en_in ? n44357_o : n44359_o;
  /* ../../HW/src/pcore/register_file.vhd:182:111  */
  assign n44359_o = dp_rd_addr[11:3];
  /* ../../HW/src/pcore/register_file.vhd:195:13  */
  assign n44364_o = wr_vector == 3'b111;
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44365_o = wr_lane[0];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44366_o = wr_lane[0];
  assign n44367_o = {n44365_o, n44366_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44368_o = wr_lane[1];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44369_o = wr_lane[1];
  assign n44370_o = {n44368_o, n44369_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44371_o = wr_lane[2];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44372_o = wr_lane[2];
  assign n44373_o = {n44371_o, n44372_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44374_o = wr_lane[3];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44375_o = wr_lane[3];
  assign n44376_o = {n44374_o, n44375_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44377_o = wr_lane[4];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44378_o = wr_lane[4];
  assign n44379_o = {n44377_o, n44378_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44380_o = wr_lane[5];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44381_o = wr_lane[5];
  assign n44382_o = {n44380_o, n44381_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44383_o = wr_lane[6];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44384_o = wr_lane[6];
  assign n44385_o = {n44383_o, n44384_o};
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44386_o = wr_lane[7];
  /* ../../HW/src/pcore/register_file.vhd:197:91  */
  assign n44387_o = wr_lane[7];
  assign n44388_o = {n44386_o, n44387_o};
  /* ../../HW/src/pcore/register_file.vhd:200:14  */
  assign n44389_o = ~wr_vector;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44391_o = 3'b000 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44392_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44393_o = n44391_o == n44392_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44396_o = n44393_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44398_o = 3'b001 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44399_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44400_o = n44398_o == n44399_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44403_o = n44400_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44405_o = 3'b010 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44406_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44407_o = n44405_o == n44406_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44410_o = n44407_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44412_o = 3'b011 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44413_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44414_o = n44412_o == n44413_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44417_o = n44414_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44419_o = 3'b100 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44420_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44421_o = n44419_o == n44420_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44424_o = n44421_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44426_o = 3'b101 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44427_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44428_o = n44426_o == n44427_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44431_o = n44428_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44433_o = 3'b110 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44434_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44435_o = n44433_o == n44434_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44438_o = n44435_o ? 2'b11 : 2'b00;
  /* ../../HW/src/pcore/register_file.vhd:202:55  */
  assign n44440_o = 3'b111 & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:77  */
  assign n44441_o = wr_vaddr & n44389_o;
  /* ../../HW/src/pcore/register_file.vhd:202:66  */
  assign n44442_o = n44440_o == n44441_o;
  /* ../../HW/src/pcore/register_file.vhd:202:4  */
  assign n44445_o = n44442_o ? 2'b11 : 2'b00;
  assign n44446_o = {n44445_o, n44438_o, n44431_o, n44424_o, n44417_o, n44410_o, n44403_o, n44396_o};
  assign n44447_o = {n44388_o, n44385_o, n44382_o, n44379_o, n44376_o, n44373_o, n44370_o, n44367_o};
  /* ../../HW/src/pcore/register_file.vhd:195:1  */
  assign n44448_o = n44364_o ? n44447_o : n44446_o;
  /* ../../HW/src/pcore/register_file.vhd:217:25  */
  assign n44454_o = wr_vector == 3'b000;
  /* ../../HW/src/pcore/register_file.vhd:218:26  */
  assign n44455_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:219:26  */
  assign n44456_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:218:56  */
  assign n44457_o = {n44455_o, n44456_o};
  /* ../../HW/src/pcore/register_file.vhd:220:26  */
  assign n44458_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:219:56  */
  assign n44459_o = {n44457_o, n44458_o};
  /* ../../HW/src/pcore/register_file.vhd:221:26  */
  assign n44460_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:220:56  */
  assign n44461_o = {n44459_o, n44460_o};
  /* ../../HW/src/pcore/register_file.vhd:222:26  */
  assign n44462_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:221:56  */
  assign n44463_o = {n44461_o, n44462_o};
  /* ../../HW/src/pcore/register_file.vhd:223:26  */
  assign n44464_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:222:56  */
  assign n44465_o = {n44463_o, n44464_o};
  /* ../../HW/src/pcore/register_file.vhd:224:26  */
  assign n44466_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:223:56  */
  assign n44467_o = {n44465_o, n44466_o};
  /* ../../HW/src/pcore/register_file.vhd:225:26  */
  assign n44468_o = wr_data[11:0];
  /* ../../HW/src/pcore/register_file.vhd:224:56  */
  assign n44469_o = {n44467_o, n44468_o};
  /* ../../HW/src/pcore/register_file.vhd:217:3  */
  assign n44470_o = n44454_o ? n44469_o : wr_data;
  /* ../../HW/src/pcore/register_file.vhd:233:16  */
  assign n44474_o = ~reset_in;
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44492_o = wr_data2[11:0];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44493_o = q1_ram_r[11:0];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44494_o = q2_ram_r[11:0];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44496_o = wr_data2[23:12];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44497_o = q1_ram_r[27:16];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44498_o = q2_ram_r[27:16];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44500_o = wr_data2[35:24];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44501_o = q1_ram_r[43:32];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44502_o = q2_ram_r[43:32];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44504_o = wr_data2[47:36];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44505_o = q1_ram_r[59:48];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44506_o = q2_ram_r[59:48];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44508_o = wr_data2[59:48];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44509_o = q1_ram_r[75:64];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44510_o = q2_ram_r[75:64];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44512_o = wr_data2[71:60];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44513_o = q1_ram_r[91:80];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44514_o = q2_ram_r[91:80];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44516_o = wr_data2[83:72];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44517_o = q1_ram_r[107:96];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44518_o = q2_ram_r[107:96];
  /* ../../HW/src/pcore/register_file.vhd:256:103  */
  assign n44520_o = wr_data2[95:84];
  /* ../../HW/src/pcore/register_file.vhd:257:85  */
  assign n44521_o = q1_ram_r[123:112];
  /* ../../HW/src/pcore/register_file.vhd:258:85  */
  assign n44522_o = q2_ram_r[123:112];
  /* ../../HW/src/pcore/register_file.vhd:264:15  */
  assign n44526_o = ~reset_in;
  /* ../../HW/src/pcore/register_file.vhd:269:10  */
  assign n44530_o = dp_read_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/register_file.vhd:343:29  */
  assign n44538_o = wr_addr[7:0];
  /* ../../HW/src/pcore/register_file.vhd:347:33  */
  assign n44539_o = rd_x1_addr[7:0];
  /* ../../HW/src/pcore/register_file.vhd:348:17  */
  assign ram3_i_n44540 = ram3_i_q1_b; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:349:33  */
  assign n44541_o = rd_x2_addr[7:0];
  /* ../../HW/src/pcore/register_file.vhd:350:17  */
  assign ram3_i_n44542 = ram3_i_q2_b; // (signal)
  /* ../../HW/src/pcore/register_file.vhd:330:1  */
  ram2r1w_256_256_8_8_128_128 ram3_i (
    .clock(clock_in),
    .clock_x2(clock_x2_in),
    .address_a(n44538_o),
    .byteena_a(byteena),
    .data_a(wr_data2_ram),
    .wren_a(wr_en),
    .address1_b(n44539_o),
    .address2_b(n44541_o),
    .q1_b(ram3_i_q1_b),
    .q2_b(ram3_i_q2_b));
  /* ../../HW/src/pcore/register_file.vhd:239:7  */
  always @(posedge clock_in or posedge n44474_o)
    if (n44474_o)
      n44547_q <= 1'b0;
    else
      n44547_q <= rd_en_in;
  /* ../../HW/src/pcore/register_file.vhd:239:7  */
  always @(posedge clock_in or posedge n44474_o)
    if (n44474_o)
      n44548_q <= 1'b0;
    else
      n44548_q <= rd_en_r;
  /* ../../HW/src/pcore/register_file.vhd:233:4  */
  assign n44549_o = {n44521_o, n44517_o, n44513_o, n44509_o, n44505_o, n44501_o, n44497_o, n44493_o};
  /* ../../HW/src/pcore/register_file.vhd:233:4  */
  assign n44550_o = {n44522_o, n44518_o, n44514_o, n44510_o, n44506_o, n44502_o, n44498_o, n44494_o};
  /* ../../HW/src/pcore/register_file.vhd:268:7  */
  always @(posedge clock_in or posedge n44526_o)
    if (n44526_o)
      n44551_q <= 1'b0;
    else
      n44551_q <= n44530_o;
  /* ../../HW/src/pcore/register_file.vhd:268:7  */
  always @(posedge clock_in or posedge n44526_o)
    if (n44526_o)
      n44552_q <= 1'b0;
    else
      n44552_q <= dp_rd_en_r;
  /* ../../HW/src/pcore/register_file.vhd:264:4  */
  assign n44553_o = {4'bX, n44520_o, 4'bX, n44516_o, 4'bX, n44512_o, 4'bX, n44508_o, 4'bX, n44504_o, 4'bX, n44500_o, 4'bX, n44496_o, 4'bX, n44492_o};
  /* ../../HW/src/pcore/register_file.vhd:239:7  */
  always @(posedge clock_in or posedge n44474_o)
    if (n44474_o)
      n44554_q <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n44554_q <= q1_ram;
  /* ../../HW/src/pcore/register_file.vhd:239:7  */
  always @(posedge clock_in or posedge n44474_o)
    if (n44474_o)
      n44555_q <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n44555_q <= q2_ram;
endmodule

module barrel_shifter_l_4_13
  (input  direction_in,
   input  [12:0] data_in,
   input  [3:0] distance_in,
   output [12:0] data_out);
  wire [3:0] distance;
  wire [12:0] shift_left;
  wire [12:0] shift_right;
  wire [12:0] n44329_o;
  wire [12:0] sra_i_n44330;
  wire [12:0] sra_i_data_out;
  wire [12:0] sla_i_n44333;
  wire [12:0] sla_i_data_out;
  assign data_out = n44329_o;
  /* ../../HW/src/util/shifter_l.vhd:42:8  */
  assign distance = distance_in; // (signal)
  /* ../../HW/src/util/shifter_l.vhd:43:8  */
  assign shift_left = sla_i_n44333; // (signal)
  /* ../../HW/src/util/shifter_l.vhd:44:8  */
  assign shift_right = sra_i_n44330; // (signal)
  /* ../../HW/src/util/shifter_l.vhd:48:25  */
  assign n44329_o = direction_in ? shift_right : shift_left;
  /* ../../HW/src/util/shifter_l.vhd:58:17  */
  assign sra_i_n44330 = sra_i_data_out; // (signal)
  /* ../../HW/src/util/shifter_l.vhd:50:1  */
  shift_right_l_4_13 sra_i (
    .data_in(data_in),
    .distance_in(distance),
    .data_out(sra_i_data_out));
  /* ../../HW/src/util/shifter_l.vhd:69:17  */
  assign sla_i_n44333 = sla_i_data_out; // (signal)
  /* ../../HW/src/util/shifter_l.vhd:61:1  */
  shift_left_l_4_13 sla_i (
    .data_in(data_in),
    .distance_in(distance),
    .data_out(sla_i_data_out));
endmodule

module barrel_shifter_a_4_13
  (input  direction_in,
   input  [12:0] data_in,
   input  [3:0] distance_in,
   output [12:0] data_out);
  wire [3:0] distance;
  wire [12:0] shift_left;
  wire [12:0] shift_right;
  wire [12:0] n44321_o;
  wire [12:0] sra_i_n44322;
  wire [12:0] sra_i_data_out;
  wire [12:0] sla_i_n44325;
  wire [12:0] sla_i_data_out;
  assign data_out = n44321_o;
  /* ../../HW/src/util/shifter.vhd:42:8  */
  assign distance = distance_in; // (signal)
  /* ../../HW/src/util/shifter.vhd:43:8  */
  assign shift_left = sla_i_n44325; // (signal)
  /* ../../HW/src/util/shifter.vhd:44:8  */
  assign shift_right = sra_i_n44322; // (signal)
  /* ../../HW/src/util/shifter.vhd:48:25  */
  assign n44321_o = direction_in ? shift_right : shift_left;
  /* ../../HW/src/util/shifter.vhd:58:17  */
  assign sra_i_n44322 = sra_i_data_out; // (signal)
  /* ../../HW/src/util/shifter.vhd:50:1  */
  shift_right_a_4_13 sra_i (
    .data_in(data_in),
    .distance_in(distance),
    .data_out(sra_i_data_out));
  /* ../../HW/src/util/shifter.vhd:69:17  */
  assign sla_i_n44325 = sla_i_data_out; // (signal)
  /* ../../HW/src/util/shifter.vhd:61:1  */
  shift_left_a_4_13 sla_i (
    .data_in(data_in),
    .distance_in(distance),
    .data_out(sla_i_data_out));
endmodule

module multiplier_13_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [12:0] x_in,
   input  [12:0] y_in,
   output [25:0] z_out);
  wire [12:0] x;
  wire [12:0] y;
  wire [25:0] z;
  wire [25:0] z_r;
  wire [25:0] n44307_o;
  wire [25:0] n44308_o;
  wire [25:0] n44309_o;
  wire n44312_o;
  wire n44317_o;
  wire [25:0] n44318_o;
  reg [25:0] n44319_q;
  assign z_out = z_r;
  /* ../../HW/src/util/multiplier.vhd:43:8  */
  assign x = x_in; // (signal)
  /* ../../HW/src/util/multiplier.vhd:44:8  */
  assign y = y_in; // (signal)
  /* ../../HW/src/util/multiplier.vhd:45:8  */
  assign z = n44309_o; // (signal)
  /* ../../HW/src/util/multiplier.vhd:46:8  */
  assign z_r = n44319_q; // (signal)
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n44307_o = {{13{x[12]}}, x}; // sext
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n44308_o = {{13{y[12]}}, y}; // sext
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n44309_o = n44307_o * n44308_o; // smul
  /* ../../HW/src/util/multiplier.vhd:63:15  */
  assign n44312_o = ~reset_in;
  /* ../../HW/src/util/multiplier.vhd:61:1  */
  assign n44317_o = ~n44312_o;
  /* ../../HW/src/util/multiplier.vhd:65:7  */
  assign n44318_o = n44317_o ? z : z_r;
  /* ../../HW/src/util/multiplier.vhd:65:7  */
  always @(posedge clock_in)
    n44319_q <= n44318_o;
endmodule

module barrel_shifter_a_2_32
  (input  direction_in,
   input  [31:0] data_in,
   input  [1:0] distance_in,
   output [31:0] data_out);
  wire [1:0] distance;
  wire [31:0] shift_left;
  wire [31:0] shift_right;
  wire [31:0] n44299_o;
  wire [31:0] sra_i_n44300;
  wire [31:0] sra_i_data_out;
  wire [31:0] sla_i_n44303;
  wire [31:0] sla_i_data_out;
  assign data_out = n44299_o;
  /* ../../HW/src/util/shifter.vhd:42:8  */
  assign distance = distance_in; // (signal)
  /* ../../HW/src/util/shifter.vhd:43:8  */
  assign shift_left = sla_i_n44303; // (signal)
  /* ../../HW/src/util/shifter.vhd:44:8  */
  assign shift_right = sra_i_n44300; // (signal)
  /* ../../HW/src/util/shifter.vhd:48:25  */
  assign n44299_o = direction_in ? shift_right : shift_left;
  /* ../../HW/src/util/shifter.vhd:58:17  */
  assign sra_i_n44300 = sra_i_data_out; // (signal)
  /* ../../HW/src/util/shifter.vhd:50:1  */
  shift_right_a_2_32 sra_i (
    .data_in(data_in),
    .distance_in(distance),
    .data_out(sra_i_data_out));
  /* ../../HW/src/util/shifter.vhd:69:17  */
  assign sla_i_n44303 = sla_i_data_out; // (signal)
  /* ../../HW/src/util/shifter.vhd:61:1  */
  shift_left_a_2_32 sla_i (
    .data_in(data_in),
    .distance_in(distance),
    .data_out(sla_i_data_out));
endmodule

module adder_32
  (input  [31:0] x_in,
   input  [31:0] y_in,
   input  add_sub_in,
   output [31:0] z_out);
  wire [31:0] x;
  wire [31:0] y;
  wire [31:0] z;
  wire [31:0] n44294_o;
  wire [31:0] n44295_o;
  wire [31:0] n44296_o;
  assign z_out = z;
  /* ../../HW/src/util/adder.vhd:38:8  */
  assign x = x_in; // (signal)
  /* ../../HW/src/util/adder.vhd:39:8  */
  assign y = y_in; // (signal)
  /* ../../HW/src/util/adder.vhd:40:8  */
  assign z = n44296_o; // (signal)
  /* ../../HW/src/util/adder.vhd:52:14  */
  assign n44294_o = x + y;
  /* ../../HW/src/util/adder.vhd:54:14  */
  assign n44295_o = x - y;
  /* ../../HW/src/util/adder.vhd:51:4  */
  assign n44296_o = add_sub_in ? n44294_o : n44295_o;
endmodule

module multiplier_12_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [11:0] x_in,
   input  [11:0] y_in,
   output [23:0] z_out);
  wire [11:0] x;
  wire [11:0] y;
  wire [23:0] z;
  wire [23:0] z_r;
  wire [23:0] n44278_o;
  wire [23:0] n44279_o;
  wire [23:0] n44280_o;
  wire n44283_o;
  wire n44288_o;
  wire [23:0] n44289_o;
  reg [23:0] n44290_q;
  assign z_out = z_r;
  /* ../../HW/src/util/multiplier.vhd:43:8  */
  assign x = x_in; // (signal)
  /* ../../HW/src/util/multiplier.vhd:44:8  */
  assign y = y_in; // (signal)
  /* ../../HW/src/util/multiplier.vhd:45:8  */
  assign z = n44280_o; // (signal)
  /* ../../HW/src/util/multiplier.vhd:46:8  */
  assign z_r = n44290_q; // (signal)
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n44278_o = {{12{x[11]}}, x}; // sext
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n44279_o = {{12{y[11]}}, y}; // sext
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n44280_o = n44278_o * n44279_o; // smul
  /* ../../HW/src/util/multiplier.vhd:63:15  */
  assign n44283_o = ~reset_in;
  /* ../../HW/src/util/multiplier.vhd:61:1  */
  assign n44288_o = ~n44283_o;
  /* ../../HW/src/util/multiplier.vhd:65:7  */
  assign n44289_o = n44288_o ? z : z_r;
  /* ../../HW/src/util/multiplier.vhd:65:7  */
  always @(posedge clock_in)
    n44290_q <= n44289_o;
endmodule

module iregister_ram_5_144
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [143:0] data1_in,
   input  [4:0] rdaddress1_in,
   input  [4:0] wraddress1_in,
   input  [17:0] wrbyteena1_in,
   input  wren1_in,
   input  rden1_in,
   output [143:0] q1_out);
  wire [143:0] data1_r;
  wire [4:0] wraddress1_r;
  wire [17:0] wrbyteena1_r;
  wire wren1_r;
  wire n44255_o;
  wire [143:0] altsyncram_i_n44270;
  wire [143:0] altsyncram_i_q_b;
  reg [143:0] n44273_q;
  reg [4:0] n44274_q;
  reg [17:0] n44275_q;
  reg n44276_q;
  assign q1_out = altsyncram_i_n44270;
  /* ../../HW/src/ialu/iregister_ram.vhd:54:8  */
  assign data1_r = n44273_q; // (signal)
  /* ../../HW/src/ialu/iregister_ram.vhd:55:8  */
  assign wraddress1_r = n44274_q; // (signal)
  /* ../../HW/src/ialu/iregister_ram.vhd:56:8  */
  assign wrbyteena1_r = n44275_q; // (signal)
  /* ../../HW/src/ialu/iregister_ram.vhd:57:8  */
  assign wren1_r = n44276_q; // (signal)
  /* ../../HW/src/ialu/iregister_ram.vhd:97:17  */
  assign n44255_o = ~reset_in;
  /* ../../HW/src/ialu/iregister_ram.vhd:127:14  */
  assign altsyncram_i_n44270 = altsyncram_i_q_b; // (signal)
  /* ../../HW/src/ialu/iregister_ram.vhd:112:1  */
  ramw_32_32_5_5_144_144 altsyncram_i (
    .clock(clock_in),
    .clock_x2(clock_x2_in),
    .address_a(wraddress1_r),
    .byteena_a(wrbyteena1_r),
    .data_a(data1_r),
    .wren_a(wren1_r),
    .address_b(rdaddress1_in),
    .q_b(altsyncram_i_q_b));
  /* ../../HW/src/ialu/iregister_ram.vhd:103:9  */
  always @(posedge clock_in or posedge n44255_o)
    if (n44255_o)
      n44273_q <= 144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n44273_q <= data1_in;
  /* ../../HW/src/ialu/iregister_ram.vhd:103:9  */
  always @(posedge clock_in or posedge n44255_o)
    if (n44255_o)
      n44274_q <= 5'b00000;
    else
      n44274_q <= wraddress1_in;
  /* ../../HW/src/ialu/iregister_ram.vhd:103:9  */
  always @(posedge clock_in or posedge n44255_o)
    if (n44255_o)
      n44275_q <= 18'b000000000000000000;
    else
      n44275_q <= wrbyteena1_in;
  /* ../../HW/src/ialu/iregister_ram.vhd:103:9  */
  always @(posedge clock_in or posedge n44255_o)
    if (n44255_o)
      n44276_q <= 1'b0;
    else
      n44276_q <= wren1_in;
endmodule

module ramw_256_256_8_8_272_272
  (input  clock,
   input  clock_x2,
   input  [7:0] address_a,
   input  [33:0] byteena_a,
   input  [271:0] data_a,
   input  wren_a,
   input  [7:0] address_b,
   output [271:0] q_b);
  wire [135:0] data;
  wire [135:0] data_r;
  wire [16:0] byteena;
  wire [16:0] byteena_r;
  wire [8:0] waddress;
  wire [7:0] waddress_r;
  wire [8:0] raddress;
  wire [7:0] raddress_r;
  wire [135:0] q;
  wire [135:0] q_latch;
  wire wren;
  wire wren_r;
  wire [135:0] n44211_o;
  wire n44212_o;
  wire [135:0] n44213_o;
  wire [16:0] n44214_o;
  wire n44215_o;
  wire [16:0] n44216_o;
  wire n44217_o;
  wire [7:0] n44218_o;
  wire n44219_o;
  wire n44220_o;
  wire [7:0] n44221_o;
  wire n44222_o;
  wire n44223_o;
  wire n44224_o;
  wire n44225_o;
  wire n44226_o;
  wire [135:0] sync_latch_i_n44227;
  wire [135:0] sync_latch_i_data_out;
  wire [135:0] n44233_o;
  wire [16:0] n44234_o;
  wire [135:0] ram_i_n44241;
  wire [135:0] ram_i_q_b;
  reg [135:0] n44244_q;
  reg [16:0] n44245_q;
  wire [8:0] n44246_o;
  reg [7:0] n44247_q;
  wire [8:0] n44248_o;
  reg [7:0] n44249_q;
  reg n44250_q;
  wire [271:0] n44251_o;
  assign q_b = n44251_o;
  /* ../../HW/src/util/ramw.vhd:55:8  */
  assign data = n44213_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:56:8  */
  assign data_r = n44244_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:57:8  */
  assign byteena = n44216_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:58:8  */
  assign byteena_r = n44245_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:59:8  */
  assign waddress = n44246_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:60:8  */
  assign waddress_r = n44247_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:61:8  */
  assign raddress = n44248_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:62:8  */
  assign raddress_r = n44249_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:63:8  */
  assign q = ram_i_n44241; // (signal)
  /* ../../HW/src/util/ramw.vhd:64:8  */
  assign q_latch = sync_latch_i_n44227; // (signal)
  /* ../../HW/src/util/ramw.vhd:65:8  */
  assign wren = n44226_o; // (signal)
  /* ../../HW/src/util/ramw.vhd:66:8  */
  assign wren_r = n44250_q; // (signal)
  /* ../../HW/src/util/ramw.vhd:69:15  */
  assign n44211_o = data_a[271:136];
  /* ../../HW/src/util/ramw.vhd:69:66  */
  assign n44212_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:69:56  */
  assign n44213_o = n44212_o ? n44211_o : data_r;
  /* ../../HW/src/util/ramw.vhd:70:21  */
  assign n44214_o = byteena_a[33:17];
  /* ../../HW/src/util/ramw.vhd:70:78  */
  assign n44215_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:70:68  */
  assign n44216_o = n44215_o ? n44214_o : byteena_r;
  /* ../../HW/src/util/ramw.vhd:71:61  */
  assign n44217_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:71:51  */
  assign n44218_o = n44217_o ? address_a : waddress_r;
  /* ../../HW/src/util/ramw.vhd:72:17  */
  assign n44219_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:73:61  */
  assign n44220_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:73:51  */
  assign n44221_o = n44220_o ? address_b : raddress_r;
  /* ../../HW/src/util/ramw.vhd:74:17  */
  assign n44222_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:77:17  */
  assign n44223_o = wren_r & clock;
  /* ../../HW/src/util/ramw.vhd:77:44  */
  assign n44224_o = ~clock;
  /* ../../HW/src/util/ramw.vhd:77:39  */
  assign n44225_o = wren_a & n44224_o;
  /* ../../HW/src/util/ramw.vhd:77:28  */
  assign n44226_o = n44223_o | n44225_o;
  /* ../../HW/src/util/ramw.vhd:88:17  */
  assign sync_latch_i_n44227 = sync_latch_i_data_out; // (signal)
  /* ../../HW/src/util/ramw.vhd:79:1  */
  sync_latch_136 sync_latch_i (
    .enable_in(clock),
    .data_in(q),
    .data_out(sync_latch_i_data_out));
  /* ../../HW/src/util/ramw.vhd:94:23  */
  assign n44233_o = data_a[135:0];
  /* ../../HW/src/util/ramw.vhd:95:29  */
  assign n44234_o = byteena_a[16:0];
  /* ../../HW/src/util/ramw.vhd:116:14  */
  assign ram_i_n44241 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/ramw.vhd:102:1  */
  dpram_be_512_512_9_9_136_136 ram_i (
    .address_a(waddress),
    .byteena_a(byteena),
    .clock0(clock_x2),
    .data_a(data),
    .wren_a(wren),
    .address_b(raddress),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n44244_q <= n44233_o;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n44245_q <= n44234_o;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  assign n44246_o = {n44218_o, n44219_o};
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n44247_q <= address_a;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  assign n44248_o = {n44221_o, n44222_o};
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n44249_q <= address_b;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  always @(posedge clock)
    n44250_q <= wren_a;
  /* ../../HW/src/util/ramw.vhd:93:4  */
  assign n44251_o = {q_latch, q};
endmodule

module dpram_512_512_9_9_132_132
  (input  [8:0] address_a,
   input  clock,
   input  [131:0] data_a,
   input  wren_a,
   input  [8:0] address_b,
   output [131:0] q_b);
  wire [8:0] address_r;
  reg [8:0] n44207_q;
  wire [131:0] n44208_data; // mem_rd
  assign q_b = n44208_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n44207_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n44207_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [131:0] ram_block[511:0] ; // memory
  assign n44208_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module dpram_256_256_8_8_67_67
  (input  [7:0] address_a,
   input  clock,
   input  [66:0] data_a,
   input  wren_a,
   input  [7:0] address_b,
   output [66:0] q_b);
  wire [7:0] address_r;
  reg [7:0] n44184_q;
  wire [66:0] n44185_data; // mem_rd
  assign q_b = n44185_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n44184_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n44184_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [66:0] ram_block[255:0] ; // memory
  assign n44185_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module dpram_32_32_5_5_388_388
  (input  [4:0] address_a,
   input  clock,
   input  [387:0] data_a,
   input  wren_a,
   input  [4:0] address_b,
   output [387:0] q_b);
  wire [4:0] address_r;
  reg [4:0] n44161_q;
  wire [387:0] n44162_data; // mem_rd
  assign q_b = n44162_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n44161_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n44161_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [387:0] ram_block[31:0] ; // memory
  assign n44162_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module sync_latch_388
  (input  enable_in,
   input  [387:0] data_in,
   output [387:0] data_out);
  wire [387:0] data_r;
  wire [387:0] n44139_o;
  assign data_out = data_r;
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:39:10  */
  assign data_r = n44139_o; // (signal)
  /* ../../HW/platform/simulation/SYNC_LATCH.vhd:45:4  */
  assign n44139_o = enable_in ? data_in : 388'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endmodule

module scfifow_1518_8
  (input  clock_in,
   input  reset_in,
   input  [1517:0] data_in,
   input  write_in,
   input  read_in,
   output writeready_out,
   output [1517:0] q_out,
   output empty_out,
   output [7:0] wused_out);
  wire [1:0] wpending_r;
  wire [1:0] rpending_r;
  wire q_avail_r;
  wire w_avail_r;
  wire [1519:0] q_r;
  wire [1519:0] data_r;
  wire [9:0] wused;
  wire write;
  wire [379:0] data;
  wire read;
  wire empty;
  wire [379:0] q;
  wire [1517:0] data_in_r;
  wire write_in_r;
  wire writeready;
  wire [379:0] fifo_i_n44014;
  wire [9:0] fifo_i_n44016;
  wire fifo_i_n44017;
  wire [379:0] fifo_i_q_out;
  wire [9:0] fifo_i_ravail_out;
  wire [9:0] fifo_i_wused_out;
  wire fifo_i_empty_out;
  wire fifo_i_full_out;
  wire fifo_i_almost_full_out;
  wire [1517:0] n44031_o;
  wire n44032_o;
  wire n44034_o;
  wire n44035_o;
  wire n44036_o;
  wire n44037_o;
  wire n44039_o;
  wire n44040_o;
  wire n44041_o;
  wire [7:0] n44042_o;
  wire [379:0] n44043_o;
  wire n44046_o;
  wire n44049_o;
  wire n44050_o;
  wire [1:0] n44052_o;
  wire n44054_o;
  wire n44056_o;
  wire [379:0] n44057_o;
  wire [379:0] n44058_o;
  wire [379:0] n44059_o;
  wire n44061_o;
  wire n44063_o;
  wire [1:0] n44065_o;
  wire [1:0] n44066_o;
  wire n44067_o;
  wire [1139:0] n44068_o;
  wire [1139:0] n44069_o;
  wire [1139:0] n44070_o;
  wire [377:0] n44071_o;
  wire [377:0] n44072_o;
  wire [377:0] n44073_o;
  wire n44074_o;
  wire n44075_o;
  wire n44076_o;
  wire [1139:0] n44077_o;
  wire n44079_o;
  wire n44081_o;
  wire [1:0] n44083_o;
  wire n44085_o;
  wire [1519:0] n44086_o;
  wire n44089_o;
  wire n44090_o;
  wire n44091_o;
  wire n44092_o;
  wire [1517:0] n44098_o;
  wire [1:0] n44116_o;
  wire [1:0] n44117_o;
  reg [1:0] n44123_q;
  wire [1:0] n44124_o;
  reg [1:0] n44125_q;
  reg n44126_q;
  reg n44127_q;
  wire [1519:0] n44128_o;
  reg [1519:0] n44129_q;
  reg [1517:0] n44130_q;
  wire [1519:0] n44131_o;
  wire [1517:0] n44132_o;
  reg [1517:0] n44133_q;
  reg n44134_q;
  assign writeready_out = writeready;
  assign q_out = n44031_o;
  assign empty_out = n44032_o;
  assign wused_out = n44042_o;
  /* ../../HW/src/util/fifow.vhd:56:8  */
  assign wpending_r = n44123_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:57:8  */
  assign rpending_r = n44125_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:58:8  */
  assign q_avail_r = n44126_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:59:8  */
  assign w_avail_r = n44127_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:60:8  */
  assign q_r = n44129_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:61:8  */
  assign data_r = n44131_o; // (signal)
  /* ../../HW/src/util/fifow.vhd:62:8  */
  assign wused = fifo_i_n44016; // (signal)
  /* ../../HW/src/util/fifow.vhd:63:8  */
  assign write = w_avail_r; // (signal)
  /* ../../HW/src/util/fifow.vhd:64:8  */
  assign data = n44043_o; // (signal)
  /* ../../HW/src/util/fifow.vhd:65:8  */
  assign read = n44037_o; // (signal)
  /* ../../HW/src/util/fifow.vhd:66:8  */
  assign empty = fifo_i_n44017; // (signal)
  /* ../../HW/src/util/fifow.vhd:67:8  */
  assign q = fifo_i_n44014; // (signal)
  /* ../../HW/src/util/fifow.vhd:70:8  */
  assign data_in_r = n44133_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:71:8  */
  assign write_in_r = n44134_q; // (signal)
  /* ../../HW/src/util/fifow.vhd:72:8  */
  assign writeready = n44041_o; // (signal)
  /* ../../HW/src/util/fifow.vhd:91:16  */
  assign fifo_i_n44014 = fifo_i_q_out; // (signal)
  /* ../../HW/src/util/fifow.vhd:93:20  */
  assign fifo_i_n44016 = fifo_i_wused_out; // (signal)
  /* ../../HW/src/util/fifow.vhd:94:20  */
  assign fifo_i_n44017 = fifo_i_empty_out; // (signal)
  /* ../../HW/src/util/fifow.vhd:76:1  */
  scfifo_380_10_4_bf8b4530d8d246dd74ac53a13471bba17941dff7 fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(data),
    .write_in(write),
    .read_in(read),
    .q_out(fifo_i_q_out),
    .ravail_out(),
    .wused_out(fifo_i_wused_out),
    .empty_out(fifo_i_empty_out),
    .full_out(),
    .almost_full_out());
  /* ../../HW/src/util/fifow.vhd:101:13  */
  assign n44031_o = q_r[1517:0];
  /* ../../HW/src/util/fifow.vhd:103:15  */
  assign n44032_o = ~q_avail_r;
  /* ../../HW/src/util/fifow.vhd:105:24  */
  assign n44034_o = ~empty;
  /* ../../HW/src/util/fifow.vhd:105:42  */
  assign n44035_o = ~q_avail_r;
  /* ../../HW/src/util/fifow.vhd:105:29  */
  assign n44036_o = n44035_o & n44034_o;
  /* ../../HW/src/util/fifow.vhd:105:13  */
  assign n44037_o = n44036_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifow.vhd:110:16  */
  assign n44039_o = ~w_avail_r;
  /* ../../HW/src/util/fifow.vhd:110:36  */
  assign n44040_o = ~write_in_r;
  /* ../../HW/src/util/fifow.vhd:110:31  */
  assign n44041_o = n44039_o & n44040_o;
  /* ../../HW/src/util/fifow.vhd:114:19  */
  assign n44042_o = wused[9:2];
  /* ../../HW/src/util/fifow.vhd:116:15  */
  assign n44043_o = data_r[379:0];
  /* ../../HW/src/util/fifow.vhd:121:15  */
  assign n44046_o = ~reset_in;
  /* ../../HW/src/util/fifow.vhd:132:10  */
  assign n44049_o = writeready ? write_in : write_in_r;
  /* ../../HW/src/util/fifow.vhd:137:22  */
  assign n44050_o = ~w_avail_r;
  /* ../../HW/src/util/fifow.vhd:139:13  */
  assign n44052_o = write_in_r ? 2'b00 : wpending_r;
  /* ../../HW/src/util/fifow.vhd:139:13  */
  assign n44054_o = write_in_r ? 1'b1 : w_avail_r;
  /* ../../HW/src/util/fifow.vhd:137:10  */
  assign n44056_o = n44074_o ? 1'b0 : n44049_o;
  /* ../../HW/src/util/fifow.vhd:146:86  */
  assign n44057_o = data_r[759:380];
  /* ../../HW/src/util/fifow.vhd:146:86  */
  assign n44058_o = data_r[1139:760];
  /* ../../HW/src/util/fifow.vhd:146:86  */
  assign n44059_o = data_r[1519:1140];
  /* ../../HW/src/util/fifow.vhd:148:26  */
  assign n44061_o = wpending_r == 2'b11;
  /* ../../HW/src/util/fifow.vhd:148:13  */
  assign n44063_o = n44061_o ? 1'b0 : w_avail_r;
  /* ../../HW/src/util/fifow.vhd:151:37  */
  assign n44065_o = wpending_r + 2'b01;
  /* ../../HW/src/util/fifow.vhd:137:10  */
  assign n44066_o = n44050_o ? n44052_o : n44065_o;
  /* ../../HW/src/util/fifow.vhd:137:10  */
  assign n44067_o = n44050_o ? n44054_o : n44063_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:285:10  */
  assign n44068_o = {n44059_o, n44058_o, n44057_o};
  assign n44069_o = data_in_r[1139:0];
  /* ../../HW/src/util/fifow.vhd:137:10  */
  assign n44070_o = n44050_o ? n44069_o : n44068_o;
  assign n44071_o = data_in_r[1517:1140];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n44072_o = data_r[1517:1140];
  /* ../../HW/src/util/fifow.vhd:137:10  */
  assign n44073_o = n44050_o ? n44071_o : n44072_o;
  /* ../../HW/src/util/fifow.vhd:137:10  */
  assign n44074_o = write_in_r & n44050_o;
  /* ../../HW/src/util/fifow.vhd:155:22  */
  assign n44075_o = ~q_avail_r;
  /* ../../HW/src/util/fifow.vhd:156:21  */
  assign n44076_o = ~empty;
  /* ../../HW/src/util/fifow.vhd:157:58  */
  assign n44077_o = q_r[1519:380];
  /* ../../HW/src/util/fifow.vhd:159:29  */
  assign n44079_o = rpending_r == 2'b11;
  /* ../../HW/src/util/fifow.vhd:156:13  */
  assign n44081_o = n44085_o ? 1'b1 : q_avail_r;
  /* ../../HW/src/util/fifow.vhd:162:40  */
  assign n44083_o = rpending_r + 2'b01;
  /* ../../HW/src/util/fifow.vhd:156:13  */
  assign n44085_o = n44079_o & n44076_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:32  */
  assign n44086_o = {q, n44077_o};
  /* ../../HW/src/util/fifow.vhd:164:10  */
  assign n44089_o = read_in ? 1'b0 : q_avail_r;
  /* ../../HW/src/util/fifow.vhd:155:10  */
  assign n44090_o = n44076_o & n44075_o;
  /* ../../HW/src/util/fifow.vhd:155:10  */
  assign n44091_o = n44075_o ? n44081_o : n44089_o;
  /* ../../HW/src/util/fifow.vhd:155:10  */
  assign n44092_o = n44076_o & n44075_o;
  assign n44098_o = {n44073_o, n44070_o};
  assign n44116_o = data_r[1519:1518];
  /* ../../HW/src/util/fifow.vhd:121:4  */
  assign n44117_o = n44046_o ? 2'b00 : n44116_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44123_q <= 2'b00;
    else
      n44123_q <= n44066_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  assign n44124_o = n44090_o ? n44083_o : rpending_r;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44125_q <= 2'b00;
    else
      n44125_q <= n44124_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44126_q <= 1'b0;
    else
      n44126_q <= n44091_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44127_q <= 1'b0;
    else
      n44127_q <= n44067_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  assign n44128_o = n44092_o ? n44086_o : q_r;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44129_q <= 1520'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n44129_q <= n44128_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44130_q <= 1518'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n44130_q <= n44098_o;
  /* ../../HW/src/util/fifow.vhd:121:4  */
  assign n44131_o = {n44117_o, n44130_q};
  /* ../../HW/src/util/fifow.vhd:131:7  */
  assign n44132_o = writeready ? data_in : data_in_r;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44133_q <= 1518'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n44133_q <= n44132_o;
  /* ../../HW/src/util/fifow.vhd:131:7  */
  always @(posedge clock_in or posedge n44046_o)
    if (n44046_o)
      n44134_q <= 1'b0;
    else
      n44134_q <= n44056_o;
endmodule

module dpram_256_256_8_8_64_64
  (input  [7:0] address_a,
   input  clock,
   input  [63:0] data_a,
   input  wren_a,
   input  [7:0] address_b,
   output [63:0] q_b);
  wire [7:0] address_r;
  reg [7:0] n44007_q;
  wire [63:0] n44008_data; // mem_rd
  assign q_b = n44008_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n44007_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n44007_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [63:0] ram_block[255:0] ; // memory
  assign n44008_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module instr_decoder2_1_3
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n42873_o;
  wire n42875_o;
  wire n42878_o;
  wire n42880_o;
  wire n42882_o;
  wire n42884_o;
  wire [5:0] n42885_o;
  wire [3:0] n42887_o;
  wire [3:0] n42889_o;
  wire [3:0] n42890_o;
  wire [3:0] n42891_o;
  reg [3:0] n42892_o;
  wire [8:0] n42894_o;
  wire [8:0] n42896_o;
  wire [8:0] n42897_o;
  wire [8:0] n42898_o;
  reg [8:0] n42899_o;
  wire [12:0] n42902_o;
  wire n42910_o;
  wire n42912_o;
  wire n42915_o;
  wire n42917_o;
  wire n42919_o;
  wire n42921_o;
  wire [5:0] n42922_o;
  wire [3:0] n42924_o;
  wire [3:0] n42926_o;
  wire [3:0] n42927_o;
  wire [3:0] n42928_o;
  reg [3:0] n42929_o;
  wire [8:0] n42931_o;
  wire [8:0] n42933_o;
  wire [8:0] n42934_o;
  wire [8:0] n42935_o;
  reg [8:0] n42936_o;
  wire [12:0] n42939_o;
  wire [7:0] n42940_o;
  wire n42941_o;
  wire [4:0] n42942_o;
  wire [4:0] n42943_o;
  wire [11:0] n42945_o;
  wire [11:0] n42946_o;
  wire [11:0] n42947_o;
  wire [11:0] n42948_o;
  wire [3:0] n42949_o;
  wire [3:0] n42950_o;
  wire [3:0] n42951_o;
  wire [3:0] n42952_o;
  wire n42953_o;
  wire n42954_o;
  wire n42955_o;
  wire n42956_o;
  wire n42959_o;
  wire n42960_o;
  wire n42961_o;
  wire n42962_o;
  wire n42963_o;
  wire n42967_o;
  wire n42968_o;
  wire n42969_o;
  wire n42970_o;
  wire n42971_o;
  wire n42975_o;
  wire n42976_o;
  wire [51:0] n42978_o;
  wire [51:0] n42979_o;
  wire [1:0] n42980_o;
  wire n42984_o;
  wire n42985_o;
  wire n42986_o;
  wire n42987_o;
  wire [12:0] n42988_o;
  wire [1:0] n42990_o;
  wire n42994_o;
  wire n42995_o;
  wire n42996_o;
  wire n42997_o;
  wire [12:0] n42998_o;
  wire [1:0] n43000_o;
  wire n43004_o;
  wire n43005_o;
  wire n43006_o;
  wire n43007_o;
  wire [12:0] n43008_o;
  wire [1:0] n43010_o;
  wire [1:0] n43014_o;
  wire [1:0] n43019_o;
  wire [1:0] n43027_o;
  wire n43031_o;
  wire n43032_o;
  wire n43033_o;
  wire n43034_o;
  wire [12:0] n43035_o;
  wire [1:0] n43037_o;
  wire n43041_o;
  wire n43042_o;
  wire [12:0] n43043_o;
  wire n43044_o;
  wire [7:0] n43045_o;
  wire [7:0] n43046_o;
  wire n43049_o;
  wire [51:0] n43051_o;
  wire [25:0] n43052_o;
  wire n43053_o;
  wire n43054_o;
  wire [12:0] n43055_o;
  wire [12:0] n43056_o;
  wire [12:0] n43057_o;
  wire n43058_o;
  wire n43059_o;
  wire [12:0] n43060_o;
  wire [12:0] n43061_o;
  wire [12:0] n43062_o;
  wire [103:0] n43073_o;
  wire [4:0] n43098_o;
  wire [3:0] n43099_o;
  wire [3:0] n43100_o;
  wire [3:0] n43101_o;
  wire [12:0] n43102_o;
  wire n43106_o;
  wire [2:0] n43108_o;
  wire [2:0] n43112_o;
  wire n43117_o;
  wire n43118_o;
  wire n43120_o;
  wire [2:0] n43121_o;
  wire [2:0] n43123_o;
  wire n43126_o;
  wire n43128_o;
  wire n43131_o;
  wire n43133_o;
  wire [2:0] n43135_o;
  wire n43137_o;
  wire n43139_o;
  wire [2:0] n43141_o;
  wire n43143_o;
  wire [4:0] n43145_o;
  wire [1:0] n43293_o;
  wire n43295_o;
  wire n43297_o;
  wire n43298_o;
  wire [2:0] n43299_o;
  wire [12:0] n43311_o;
  wire [12:0] n43312_o;
  wire [12:0] n43313_o;
  wire [9:0] n43315_o;
  wire [12:0] n43319_o;
  wire [12:0] n43320_o;
  wire [12:0] n43322_o;
  wire [9:0] n43324_o;
  wire [12:0] n43328_o;
  wire [12:0] n43329_o;
  wire n43331_o;
  wire [1:0] n43332_o;
  wire n43334_o;
  wire n43335_o;
  wire [11:0] n43336_o;
  wire [8:0] n43337_o;
  wire [8:0] n43338_o;
  wire [2:0] n43339_o;
  wire [2:0] n43340_o;
  wire [2:0] n43341_o;
  wire n43343_o;
  wire [1:0] n43344_o;
  wire n43346_o;
  wire n43347_o;
  wire n43349_o;
  wire n43350_o;
  wire n43352_o;
  wire [4:0] n43353_o;
  wire [8:0] n43354_o;
  wire [4:0] n43355_o;
  wire [5:0] n43357_o;
  wire [2:0] n43358_o;
  wire [8:0] n43359_o;
  wire [8:0] n43360_o;
  wire [2:0] n43361_o;
  wire [12:0] n43362_o;
  wire n43363_o;
  wire [11:0] n43364_o;
  wire [8:0] n43365_o;
  wire [8:0] n43366_o;
  wire [2:0] n43367_o;
  wire n43369_o;
  wire [4:0] n43370_o;
  wire [8:0] n43371_o;
  wire [4:0] n43372_o;
  wire [5:0] n43374_o;
  wire [2:0] n43375_o;
  wire [8:0] n43376_o;
  wire [8:0] n43377_o;
  wire [2:0] n43378_o;
  wire [11:0] n43379_o;
  wire [11:0] n43380_o;
  wire [11:0] n43381_o;
  wire [11:0] n43382_o;
  wire [11:0] n43383_o;
  wire [11:0] n43386_o;
  wire [11:0] n43387_o;
  wire [1:0] n43403_o;
  wire n43405_o;
  wire n43407_o;
  wire n43408_o;
  wire [2:0] n43409_o;
  wire [12:0] n43421_o;
  wire [12:0] n43422_o;
  wire [12:0] n43423_o;
  wire [9:0] n43425_o;
  wire [12:0] n43429_o;
  wire [12:0] n43430_o;
  wire [12:0] n43432_o;
  wire [9:0] n43434_o;
  wire [12:0] n43438_o;
  wire [12:0] n43439_o;
  wire n43441_o;
  wire [1:0] n43442_o;
  wire n43444_o;
  wire n43445_o;
  wire [11:0] n43446_o;
  wire [8:0] n43447_o;
  wire [8:0] n43448_o;
  wire [2:0] n43449_o;
  wire [2:0] n43450_o;
  wire [2:0] n43451_o;
  wire n43453_o;
  wire [1:0] n43454_o;
  wire n43456_o;
  wire n43457_o;
  wire n43459_o;
  wire n43460_o;
  wire n43462_o;
  wire [4:0] n43463_o;
  wire [8:0] n43464_o;
  wire [4:0] n43465_o;
  wire [5:0] n43467_o;
  wire [2:0] n43468_o;
  wire [8:0] n43469_o;
  wire [8:0] n43470_o;
  wire [2:0] n43471_o;
  wire [12:0] n43472_o;
  wire n43473_o;
  wire [11:0] n43474_o;
  wire [8:0] n43475_o;
  wire [8:0] n43476_o;
  wire [2:0] n43477_o;
  wire n43479_o;
  wire [4:0] n43480_o;
  wire [8:0] n43481_o;
  wire [4:0] n43482_o;
  wire [5:0] n43484_o;
  wire [2:0] n43485_o;
  wire [8:0] n43486_o;
  wire [8:0] n43487_o;
  wire [2:0] n43488_o;
  wire [11:0] n43489_o;
  wire [11:0] n43490_o;
  wire [11:0] n43491_o;
  wire [11:0] n43492_o;
  wire [11:0] n43493_o;
  wire [11:0] n43496_o;
  wire [11:0] n43497_o;
  wire [1:0] n43513_o;
  wire n43515_o;
  wire n43517_o;
  wire n43518_o;
  wire [2:0] n43519_o;
  wire [12:0] n43531_o;
  wire [12:0] n43532_o;
  wire [12:0] n43533_o;
  wire [9:0] n43535_o;
  wire [12:0] n43539_o;
  wire [12:0] n43540_o;
  wire [12:0] n43542_o;
  wire [9:0] n43544_o;
  wire [12:0] n43548_o;
  wire [12:0] n43549_o;
  wire n43551_o;
  wire [1:0] n43552_o;
  wire n43554_o;
  wire n43555_o;
  wire [11:0] n43556_o;
  wire [8:0] n43557_o;
  wire [8:0] n43558_o;
  wire [2:0] n43559_o;
  wire [2:0] n43560_o;
  wire [2:0] n43561_o;
  wire n43563_o;
  wire [1:0] n43564_o;
  wire n43566_o;
  wire n43567_o;
  wire n43569_o;
  wire n43570_o;
  wire n43572_o;
  wire [4:0] n43573_o;
  wire [8:0] n43574_o;
  wire [4:0] n43575_o;
  wire [5:0] n43577_o;
  wire [2:0] n43578_o;
  wire [8:0] n43579_o;
  wire [8:0] n43580_o;
  wire [2:0] n43581_o;
  wire [12:0] n43582_o;
  wire n43583_o;
  wire [11:0] n43584_o;
  wire [8:0] n43585_o;
  wire [8:0] n43586_o;
  wire [2:0] n43587_o;
  wire n43589_o;
  wire [4:0] n43590_o;
  wire [8:0] n43591_o;
  wire [4:0] n43592_o;
  wire [5:0] n43594_o;
  wire [2:0] n43595_o;
  wire [8:0] n43596_o;
  wire [8:0] n43597_o;
  wire [2:0] n43598_o;
  wire [11:0] n43599_o;
  wire [11:0] n43600_o;
  wire [11:0] n43601_o;
  wire [11:0] n43602_o;
  wire [11:0] n43603_o;
  wire [11:0] n43606_o;
  wire [11:0] n43607_o;
  wire [1:0] n43623_o;
  wire n43625_o;
  wire n43627_o;
  wire n43628_o;
  wire [2:0] n43629_o;
  wire [12:0] n43641_o;
  wire [12:0] n43642_o;
  wire [12:0] n43643_o;
  wire [9:0] n43645_o;
  wire [12:0] n43649_o;
  wire [12:0] n43650_o;
  wire [12:0] n43652_o;
  wire [9:0] n43654_o;
  wire [12:0] n43658_o;
  wire [12:0] n43659_o;
  wire n43661_o;
  wire [1:0] n43662_o;
  wire n43664_o;
  wire n43665_o;
  wire [11:0] n43666_o;
  wire [8:0] n43667_o;
  wire [8:0] n43668_o;
  wire [2:0] n43669_o;
  wire [2:0] n43670_o;
  wire [2:0] n43671_o;
  wire n43673_o;
  wire [1:0] n43674_o;
  wire n43676_o;
  wire n43677_o;
  wire n43679_o;
  wire n43680_o;
  wire n43682_o;
  wire [4:0] n43683_o;
  wire [8:0] n43684_o;
  wire [4:0] n43685_o;
  wire [5:0] n43687_o;
  wire [2:0] n43688_o;
  wire [8:0] n43689_o;
  wire [8:0] n43690_o;
  wire [2:0] n43691_o;
  wire [12:0] n43692_o;
  wire n43693_o;
  wire [11:0] n43694_o;
  wire [8:0] n43695_o;
  wire [8:0] n43696_o;
  wire [2:0] n43697_o;
  wire n43699_o;
  wire [4:0] n43700_o;
  wire [8:0] n43701_o;
  wire [4:0] n43702_o;
  wire [5:0] n43704_o;
  wire [2:0] n43705_o;
  wire [8:0] n43706_o;
  wire [8:0] n43707_o;
  wire [2:0] n43708_o;
  wire [11:0] n43709_o;
  wire [11:0] n43710_o;
  wire [11:0] n43711_o;
  wire [11:0] n43712_o;
  wire [11:0] n43713_o;
  wire [11:0] n43716_o;
  wire [11:0] n43717_o;
  wire n43724_o;
  wire [11:0] n43726_o;
  wire [6:0] n43727_o;
  wire [7:0] n43728_o;
  wire [3:0] n43730_o;
  wire [7:0] n43731_o;
  wire [6:0] n43732_o;
  wire [7:0] n43733_o;
  wire [7:0] n43734_o;
  wire n43737_o;
  wire n43739_o;
  wire n43741_o;
  wire n43743_o;
  wire n43745_o;
  wire [4:0] n43747_o;
  wire [7:0] n43752_o;
  wire [7:0] n43754_o;
  wire [7:0] n43756_o;
  wire [7:0] n43758_o;
  reg [3:0] n43829_q;
  reg [3:0] n43830_q;
  reg [3:0] n43831_q;
  reg [3:0] n43832_q;
  reg [3:0] n43833_q;
  reg [3:0] n43834_q;
  reg n43836_q;
  reg n43837_q;
  reg [12:0] n43838_q;
  reg [12:0] n43839_q;
  reg [12:0] n43840_q;
  reg n43841_q;
  reg n43842_q;
  reg n43843_q;
  reg n43844_q;
  reg n43846_q;
  reg n43847_q;
  reg n43848_q;
  reg n43849_q;
  reg n43850_q;
  reg n43851_q;
  reg [11:0] n43852_q;
  reg n43853_q;
  reg n43854_q;
  reg n43855_q;
  reg [4:0] n43856_q;
  wire [11:0] n43857_o;
  reg [11:0] n43858_q;
  wire [11:0] n43859_o;
  reg [11:0] n43860_q;
  wire [11:0] n43861_o;
  reg [11:0] n43862_q;
  reg n43863_q;
  reg n43864_q;
  reg n43865_q;
  reg n43866_q;
  reg n43867_q;
  reg n43868_q;
  reg [4:0] n43870_q;
  reg [3:0] n43871_q;
  reg [3:0] n43872_q;
  reg [3:0] n43873_q;
  reg [12:0] n43874_q;
  reg [4:0] n43875_q;
  reg [3:0] n43876_q;
  reg [3:0] n43877_q;
  reg [3:0] n43878_q;
  reg [3:0] n43879_q;
  reg [3:0] n43880_q;
  reg [12:0] n43881_q;
  reg [12:0] n43882_q;
  reg [2:0] n43883_q;
  reg [2:0] n43884_q;
  reg [2:0] n43885_q;
  reg [2:0] n43886_q;
  reg n43888_q;
  reg n43889_q;
  reg n43890_q;
  reg n43891_q;
  reg [4:0] n43893_q;
  reg [103:0] n43894_q;
  reg [12:0] n43895_q;
  reg [12:0] n43896_q;
  reg [12:0] n43897_q;
  reg [12:0] n43898_q;
  reg [12:0] n43899_q;
  reg [12:0] n43900_q;
  reg [7:0] n43901_q;
  reg [7:0] n43902_q;
  reg [7:0] n43903_q;
  reg [7:0] n43904_q;
  reg [7:0] n43905_q;
  reg [7:0] n43906_q;
  reg [7:0] n43907_q;
  reg [7:0] n43908_q;
  reg [7:0] n43909_q;
  reg [12:0] n43910_q;
  wire [12:0] n43911_o;
  wire [12:0] n43912_o;
  wire [12:0] n43913_o;
  wire [12:0] n43914_o;
  wire [1:0] n43915_o;
  reg [12:0] n43916_o;
  wire [12:0] n43917_o;
  wire [12:0] n43918_o;
  wire [12:0] n43919_o;
  wire [12:0] n43920_o;
  wire [1:0] n43921_o;
  reg [12:0] n43922_o;
  wire [12:0] n43923_o;
  wire [12:0] n43924_o;
  wire [12:0] n43925_o;
  wire [12:0] n43926_o;
  wire [1:0] n43927_o;
  reg [12:0] n43928_o;
  wire [12:0] n43929_o;
  wire [12:0] n43930_o;
  wire [12:0] n43931_o;
  wire [12:0] n43932_o;
  wire [1:0] n43933_o;
  reg [12:0] n43934_o;
  wire [12:0] n43935_o;
  wire [12:0] n43936_o;
  wire [12:0] n43937_o;
  wire [12:0] n43938_o;
  wire [1:0] n43939_o;
  reg [12:0] n43940_o;
  wire [12:0] n43941_o;
  wire [12:0] n43942_o;
  wire [12:0] n43943_o;
  wire [12:0] n43944_o;
  wire [1:0] n43945_o;
  reg [12:0] n43946_o;
  wire [12:0] n43947_o;
  wire [12:0] n43948_o;
  wire [12:0] n43949_o;
  wire [12:0] n43950_o;
  wire [1:0] n43951_o;
  reg [12:0] n43952_o;
  wire [12:0] n43953_o;
  wire [12:0] n43954_o;
  wire [12:0] n43955_o;
  wire [12:0] n43956_o;
  wire [1:0] n43957_o;
  reg [12:0] n43958_o;
  wire [12:0] n43959_o;
  wire [12:0] n43960_o;
  wire [12:0] n43961_o;
  wire [12:0] n43962_o;
  wire [12:0] n43963_o;
  wire [12:0] n43964_o;
  wire [12:0] n43965_o;
  wire [12:0] n43966_o;
  wire [1:0] n43967_o;
  reg [12:0] n43968_o;
  wire [1:0] n43969_o;
  reg [12:0] n43970_o;
  wire n43971_o;
  wire [12:0] n43972_o;
  wire [12:0] n43973_o;
  wire [12:0] n43974_o;
  wire [12:0] n43975_o;
  wire [12:0] n43976_o;
  wire [12:0] n43977_o;
  wire [12:0] n43978_o;
  wire [12:0] n43979_o;
  wire [12:0] n43980_o;
  wire [1:0] n43981_o;
  reg [12:0] n43982_o;
  wire [1:0] n43983_o;
  reg [12:0] n43984_o;
  wire n43985_o;
  wire [12:0] n43986_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n43045_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n42902_o;
  assign i_x2_out = n42939_o;
  assign result_waddr_out = n42940_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n43829_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n43830_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n43831_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n43832_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n43833_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n43834_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n43836_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n43837_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n43838_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n43839_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n43840_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n43841_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n43842_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n43843_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n43844_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n42943_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n43846_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n43847_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n42941_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n43848_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n42963_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n43849_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n42971_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n43850_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n42976_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n43851_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n43852_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n42945_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n42946_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n42947_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n42948_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n42949_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n42950_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n42951_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n42952_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n42953_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n42954_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n42955_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n42956_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n43853_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n43854_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n43855_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n43856_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n43858_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n43860_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n43862_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n43387_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n43497_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n43607_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n43717_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n43863_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n43864_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n43865_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n43866_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n43867_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n43868_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n43098_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n43099_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n43100_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n43101_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n43102_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n43870_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n43871_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n43872_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n43873_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n43874_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n43875_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n43876_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n43877_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n43878_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n43879_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n43880_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n43881_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n43882_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n43883_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n43884_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n43885_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n43886_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n43888_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n43889_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n43890_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n43891_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n43893_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n43894_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n42978_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n42979_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n43895_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n43896_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n43897_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n43898_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n43899_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n43900_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n42988_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n42998_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n43008_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n43934_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n43940_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n43946_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n43043_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n43035_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n43958_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n43901_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n43902_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n43903_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n43904_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n43905_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n43906_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n43907_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n43908_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n43909_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n43910_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n42873_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n42875_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n42878_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n42880_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n42882_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n42884_o = imu_x1_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42885_o = {n42884_o, n42882_o, n42880_o, n42878_o, n42875_o, n42873_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42887_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42889_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42890_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42891_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n42885_o)
      6'b100000: n42892_o = n42890_o;
      6'b010000: n42892_o = n42889_o;
      6'b001000: n42892_o = 4'b0111;
      6'b000100: n42892_o = instruction_tid_rrr;
      6'b000010: n42892_o = n42887_o;
      6'b000001: n42892_o = 4'b0000;
      default: n42892_o = n42891_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42894_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42896_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42897_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42898_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n42885_o)
      6'b100000: n42899_o = n42897_o;
      6'b010000: n42899_o = n42896_o;
      6'b001000: n42899_o = 9'b000000000;
      6'b000100: n42899_o = 9'b000000000;
      6'b000010: n42899_o = n42894_o;
      6'b000001: n42899_o = 9'b000000000;
      default: n42899_o = n42898_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42902_o = {n42899_o, n42892_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n42910_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n42912_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n42915_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n42917_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n42919_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n42921_o = imu_x2_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42922_o = {n42921_o, n42919_o, n42917_o, n42915_o, n42912_o, n42910_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42924_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42926_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42927_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n42928_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n42922_o)
      6'b100000: n42929_o = n42927_o;
      6'b010000: n42929_o = n42926_o;
      6'b001000: n42929_o = 4'b0111;
      6'b000100: n42929_o = instruction_tid_rrr;
      6'b000010: n42929_o = n42924_o;
      6'b000001: n42929_o = 4'b0000;
      default: n42929_o = n42928_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42931_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42933_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42934_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42935_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n42922_o)
      6'b100000: n42936_o = n42934_o;
      6'b010000: n42936_o = n42933_o;
      6'b001000: n42936_o = 9'b000000000;
      6'b000100: n42936_o = 9'b000000000;
      6'b000010: n42936_o = n42931_o;
      6'b000001: n42936_o = 9'b000000000;
      default: n42936_o = n42935_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n42939_o = {n42936_o, n42929_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n42940_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n42941_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n42942_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n42943_o = instruction_mu_valid_in ? n42942_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n42945_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n42946_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n42947_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n42948_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n42949_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n42950_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n42951_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n42952_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n42953_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n42954_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n42955_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n42956_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n42959_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n42960_o = n42959_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n42961_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n42962_o = n42961_o & n42960_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n42963_o = n42962_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n42967_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n42968_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n42969_o = n42968_o & n42967_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n42970_o = n42969_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n42971_o = n42970_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n42975_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n42976_o = n42975_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n42978_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n42979_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n42980_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n42984_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n42985_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n42986_o = ~n42985_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n42987_o = n42984_o | n42986_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n42988_o = n42987_o ? n43916_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n42990_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n42994_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n42995_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n42996_o = ~n42995_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n42997_o = n42994_o | n42996_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n42998_o = n42997_o ? n43922_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n43000_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n43004_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n43005_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n43006_o = ~n43005_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n43007_o = n43004_o | n43006_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n43008_o = n43007_o ? n43928_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n43010_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n43014_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n43019_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n43027_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n43031_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n43032_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n43033_o = ~n43032_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n43034_o = n43031_o | n43033_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n43035_o = n43034_o ? n43952_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n43037_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n43041_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n43042_o = ~n43041_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n43043_o = n43042_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n43044_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n43045_o = n43044_o ? mu_lane_rrrrrr : n43046_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n43046_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n43049_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n43051_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n43052_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n43053_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n43054_o = ~n43053_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n43055_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n43056_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n43057_o = n43054_o ? n43055_o : n43056_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n43058_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n43059_o = ~n43058_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n43060_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n43061_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n43062_o = n43059_o ? n43060_o : n43061_o;
  assign n43073_o = {n43051_o, n43057_o, n43062_o, n43052_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n43098_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n43099_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n43100_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n43101_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n43102_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n43106_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n43108_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n43112_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n43117_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n43118_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n43120_o = n43118_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n43121_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n43123_o = n43120_o ? n43121_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n43126_o = n43120_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n43128_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n43131_o = n43128_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n43133_o = n43117_o ? n43131_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n43135_o = n43117_o ? n43123_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n43137_o = n43117_o ? n43126_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n43139_o = got_imu_rr ? n43133_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n43141_o = got_imu_rr ? n43135_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n43143_o = got_imu_rr ? n43137_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n43145_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n43293_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n43295_o = n43293_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n43297_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n43298_o = n43295_o | n43297_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n43299_o = mu_x1_parm1[2:0];
  assign n43311_o = {1'b0, mu_x1_parm1};
  assign n43312_o = {10'b0000000000, n43299_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n43313_o = n43298_o ? n43312_o : n43311_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n43315_o = mu_x1_i1_1[9:0];
  assign n43319_o = {n43315_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n43320_o = mu_x1_vector ? n43319_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n43322_o = mu_x1_i0_1 + n43313_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n43324_o = n43322_o[9:0];
  assign n43328_o = {n43324_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43329_o = mu_x1_vector ? n43328_o : n43322_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n43331_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n43332_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n43334_o = n43332_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n43335_o = n43331_o | n43334_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n43336_o = n43329_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n43337_o = n43336_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n43338_o = ~n43337_o;
  assign n43339_o = n43328_o[2:0];
  assign n43340_o = n43322_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43341_o = mu_x1_vector ? n43339_o : n43340_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n43343_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n43344_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n43346_o = n43344_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n43347_o = n43343_o | n43346_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n43349_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n43350_o = n43347_o | n43349_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n43352_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n43353_o = n43329_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n43354_o = {n43353_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n43355_o = n43329_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n43357_o = {1'b0, n43355_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n43358_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n43359_o = {n43357_o, n43358_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n43360_o = n43352_o ? n43354_o : n43359_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n43361_o = n43329_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n43362_o = n43320_o + n43329_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n43363_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n43364_o = n43362_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n43365_o = n43364_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n43366_o = ~n43365_o;
  assign n43367_o = n43362_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n43369_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n43370_o = n43362_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n43371_o = {n43370_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n43372_o = n43362_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n43374_o = {1'b0, n43372_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n43375_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n43376_o = {n43374_o, n43375_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n43377_o = n43369_o ? n43371_o : n43376_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n43378_o = n43362_o[2:0];
  assign n43379_o = {n43377_o, n43378_o};
  assign n43380_o = {n43366_o, n43367_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n43381_o = n43363_o ? n43380_o : n43379_o;
  assign n43382_o = {n43360_o, n43361_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n43383_o = n43350_o ? n43382_o : n43381_o;
  assign n43386_o = {n43338_o, n43341_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n43387_o = n43335_o ? n43386_o : n43383_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n43403_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n43405_o = n43403_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n43407_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n43408_o = n43405_o | n43407_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n43409_o = mu_x2_parm1[2:0];
  assign n43421_o = {1'b0, mu_x2_parm1};
  assign n43422_o = {10'b0000000000, n43409_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n43423_o = n43408_o ? n43422_o : n43421_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n43425_o = mu_x2_i1_1[9:0];
  assign n43429_o = {n43425_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n43430_o = mu_x2_vector ? n43429_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n43432_o = mu_x2_i0_1 + n43423_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n43434_o = n43432_o[9:0];
  assign n43438_o = {n43434_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43439_o = mu_x2_vector ? n43438_o : n43432_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n43441_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n43442_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n43444_o = n43442_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n43445_o = n43441_o | n43444_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n43446_o = n43439_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n43447_o = n43446_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n43448_o = ~n43447_o;
  assign n43449_o = n43438_o[2:0];
  assign n43450_o = n43432_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43451_o = mu_x2_vector ? n43449_o : n43450_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n43453_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n43454_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n43456_o = n43454_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n43457_o = n43453_o | n43456_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n43459_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n43460_o = n43457_o | n43459_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n43462_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n43463_o = n43439_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n43464_o = {n43463_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n43465_o = n43439_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n43467_o = {1'b0, n43465_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n43468_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n43469_o = {n43467_o, n43468_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n43470_o = n43462_o ? n43464_o : n43469_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n43471_o = n43439_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n43472_o = n43430_o + n43439_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n43473_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n43474_o = n43472_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n43475_o = n43474_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n43476_o = ~n43475_o;
  assign n43477_o = n43472_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n43479_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n43480_o = n43472_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n43481_o = {n43480_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n43482_o = n43472_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n43484_o = {1'b0, n43482_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n43485_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n43486_o = {n43484_o, n43485_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n43487_o = n43479_o ? n43481_o : n43486_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n43488_o = n43472_o[2:0];
  assign n43489_o = {n43487_o, n43488_o};
  assign n43490_o = {n43476_o, n43477_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n43491_o = n43473_o ? n43490_o : n43489_o;
  assign n43492_o = {n43470_o, n43471_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n43493_o = n43460_o ? n43492_o : n43491_o;
  assign n43496_o = {n43448_o, n43451_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n43497_o = n43445_o ? n43496_o : n43493_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n43513_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n43515_o = n43513_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n43517_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n43518_o = n43515_o | n43517_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n43519_o = mu_x3_parm1[2:0];
  assign n43531_o = {1'b0, mu_x3_parm1};
  assign n43532_o = {10'b0000000000, n43519_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n43533_o = n43518_o ? n43532_o : n43531_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n43535_o = mu_x3_i1_1[9:0];
  assign n43539_o = {n43535_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n43540_o = mu_x3_vector ? n43539_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n43542_o = mu_x3_i0_1 + n43533_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n43544_o = n43542_o[9:0];
  assign n43548_o = {n43544_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43549_o = mu_x3_vector ? n43548_o : n43542_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n43551_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n43552_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n43554_o = n43552_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n43555_o = n43551_o | n43554_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n43556_o = n43549_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n43557_o = n43556_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n43558_o = ~n43557_o;
  assign n43559_o = n43548_o[2:0];
  assign n43560_o = n43542_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43561_o = mu_x3_vector ? n43559_o : n43560_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n43563_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n43564_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n43566_o = n43564_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n43567_o = n43563_o | n43566_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n43569_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n43570_o = n43567_o | n43569_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n43572_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n43573_o = n43549_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n43574_o = {n43573_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n43575_o = n43549_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n43577_o = {1'b0, n43575_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n43578_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n43579_o = {n43577_o, n43578_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n43580_o = n43572_o ? n43574_o : n43579_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n43581_o = n43549_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n43582_o = n43540_o + n43549_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n43583_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n43584_o = n43582_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n43585_o = n43584_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n43586_o = ~n43585_o;
  assign n43587_o = n43582_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n43589_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n43590_o = n43582_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n43591_o = {n43590_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n43592_o = n43582_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n43594_o = {1'b0, n43592_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n43595_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n43596_o = {n43594_o, n43595_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n43597_o = n43589_o ? n43591_o : n43596_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n43598_o = n43582_o[2:0];
  assign n43599_o = {n43597_o, n43598_o};
  assign n43600_o = {n43586_o, n43587_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n43601_o = n43583_o ? n43600_o : n43599_o;
  assign n43602_o = {n43580_o, n43581_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n43603_o = n43570_o ? n43602_o : n43601_o;
  assign n43606_o = {n43558_o, n43561_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n43607_o = n43555_o ? n43606_o : n43603_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n43623_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n43625_o = n43623_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n43627_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n43628_o = n43625_o | n43627_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n43629_o = mu_y_parm1[2:0];
  assign n43641_o = {1'b0, mu_y_parm1};
  assign n43642_o = {10'b0000000000, n43629_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n43643_o = n43628_o ? n43642_o : n43641_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n43645_o = mu_y_i1_1[9:0];
  assign n43649_o = {n43645_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n43650_o = mu_y_vector ? n43649_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n43652_o = mu_y_i0_1 + n43643_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n43654_o = n43652_o[9:0];
  assign n43658_o = {n43654_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43659_o = mu_y_vector ? n43658_o : n43652_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n43661_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n43662_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n43664_o = n43662_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n43665_o = n43661_o | n43664_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n43666_o = n43659_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n43667_o = n43666_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n43668_o = ~n43667_o;
  assign n43669_o = n43658_o[2:0];
  assign n43670_o = n43652_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n43671_o = mu_y_vector ? n43669_o : n43670_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n43673_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n43674_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n43676_o = n43674_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n43677_o = n43673_o | n43676_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n43679_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n43680_o = n43677_o | n43679_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n43682_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n43683_o = n43659_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n43684_o = {n43683_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n43685_o = n43659_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n43687_o = {1'b0, n43685_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n43688_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n43689_o = {n43687_o, n43688_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n43690_o = n43682_o ? n43684_o : n43689_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n43691_o = n43659_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n43692_o = n43650_o + n43659_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n43693_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n43694_o = n43692_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n43695_o = n43694_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n43696_o = ~n43695_o;
  assign n43697_o = n43692_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n43699_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n43700_o = n43692_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n43701_o = {n43700_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n43702_o = n43692_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n43704_o = {1'b0, n43702_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n43705_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n43706_o = {n43704_o, n43705_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n43707_o = n43699_o ? n43701_o : n43706_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n43708_o = n43692_o[2:0];
  assign n43709_o = {n43707_o, n43708_o};
  assign n43710_o = {n43696_o, n43697_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n43711_o = n43693_o ? n43710_o : n43709_o;
  assign n43712_o = {n43690_o, n43691_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n43713_o = n43680_o ? n43712_o : n43711_o;
  assign n43716_o = {n43668_o, n43671_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n43717_o = n43665_o ? n43716_o : n43713_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n43724_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n43726_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n43727_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n43728_o = {instruction_vm_in, n43727_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n43730_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n43731_o = {n43730_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n43732_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n43733_o = {instruction_vm_in, n43732_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n43734_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43737_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43739_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43741_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43743_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43745_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43747_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43752_o = instruction_tid_valid_in ? n43734_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43754_o = instruction_tid_valid_in ? n43733_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43756_o = instruction_tid_valid_in ? n43731_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n43758_o = instruction_tid_valid_in ? n43728_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43829_q <= 4'b0000;
    else
      n43829_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43830_q <= 4'b0000;
    else
      n43830_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43831_q <= 4'b0000;
    else
      n43831_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43832_q <= 4'b0000;
    else
      n43832_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43833_q <= 4'b0000;
    else
      n43833_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43834_q <= 4'b0000;
    else
      n43834_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43836_q <= 1'b0;
    else
      n43836_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43837_q <= 1'b0;
    else
      n43837_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43838_q <= 13'b0000000000000;
    else
      n43838_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43839_q <= 13'b0000000000000;
    else
      n43839_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43840_q <= 13'b0000000000000;
    else
      n43840_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43841_q <= 1'b0;
    else
      n43841_q <= n43139_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43842_q <= 1'b0;
    else
      n43842_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43843_q <= 1'b0;
    else
      n43843_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43844_q <= 1'b0;
    else
      n43844_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43846_q <= 1'b0;
    else
      n43846_q <= n43737_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43847_q <= 1'b0;
    else
      n43847_q <= n43739_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43848_q <= 1'b0;
    else
      n43848_q <= n43741_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43849_q <= 1'b0;
    else
      n43849_q <= n43743_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43850_q <= 1'b0;
    else
      n43850_q <= n43745_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43851_q <= 1'b0;
    else
      n43851_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43852_q <= 12'b000000000000;
    else
      n43852_q <= n43726_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43853_q <= 1'b0;
    else
      n43853_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43854_q <= 1'b0;
    else
      n43854_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43855_q <= 1'b0;
    else
      n43855_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43856_q <= 5'b00000;
    else
      n43856_q <= n43747_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n43857_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43858_q <= 12'b000000000000;
    else
      n43858_q <= n43857_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n43859_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43860_q <= 12'b000000000000;
    else
      n43860_q <= n43859_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n43861_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43862_q <= 12'b000000000000;
    else
      n43862_q <= n43861_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43863_q <= 1'b0;
    else
      n43863_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43864_q <= 1'b0;
    else
      n43864_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43865_q <= 1'b0;
    else
      n43865_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43866_q <= 1'b0;
    else
      n43866_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43867_q <= 1'b0;
    else
      n43867_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43868_q <= 1'b0;
    else
      n43868_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43870_q <= 5'b00000;
    else
      n43870_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43871_q <= 4'b0000;
    else
      n43871_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43872_q <= 4'b0000;
    else
      n43872_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43873_q <= 4'b0000;
    else
      n43873_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43874_q <= 13'b0000000000000;
    else
      n43874_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43875_q <= 5'b00000;
    else
      n43875_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43876_q <= 4'b0000;
    else
      n43876_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43877_q <= 4'b0000;
    else
      n43877_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43878_q <= 4'b0000;
    else
      n43878_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43879_q <= 4'b0000;
    else
      n43879_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43880_q <= 4'b0000;
    else
      n43880_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43881_q <= 13'b0000000000000;
    else
      n43881_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43882_q <= 13'b0000000000000;
    else
      n43882_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43883_q <= 3'b000;
    else
      n43883_q <= n43141_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43884_q <= 3'b000;
    else
      n43884_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43885_q <= 3'b000;
    else
      n43885_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43886_q <= 3'b000;
    else
      n43886_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43888_q <= 1'b0;
    else
      n43888_q <= n43143_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43889_q <= 1'b0;
    else
      n43889_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43890_q <= 1'b0;
    else
      n43890_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43891_q <= 1'b0;
    else
      n43891_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43893_q <= 5'b00000;
    else
      n43893_q <= n43145_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n43049_o)
    if (n43049_o)
      n43894_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n43894_q <= n43073_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43895_q <= 13'b0000000000000;
    else
      n43895_q <= n43972_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43896_q <= 13'b0000000000000;
    else
      n43896_q <= n43986_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43897_q <= 13'b0000000000000;
    else
      n43897_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43898_q <= 13'b0000000000000;
    else
      n43898_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43899_q <= 13'b0000000000000;
    else
      n43899_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43900_q <= 13'b0000000000000;
    else
      n43900_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43901_q <= 8'b00000000;
    else
      n43901_q <= n43752_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43902_q <= 8'b00000000;
    else
      n43902_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43903_q <= 8'b00000000;
    else
      n43903_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43904_q <= 8'b00000000;
    else
      n43904_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43905_q <= 8'b00000000;
    else
      n43905_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43906_q <= 8'b00000000;
    else
      n43906_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43907_q <= 8'b00000000;
    else
      n43907_q <= n43754_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43908_q <= 8'b00000000;
    else
      n43908_q <= n43756_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n43724_o)
    if (n43724_o)
      n43909_q <= 8'b00000000;
    else
      n43909_q <= n43758_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n43106_o)
    if (n43106_o)
      n43910_q <= 13'b0000000000000;
    else
      n43910_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n43911_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n43912_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n43913_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n43914_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n43915_o = n42980_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n43915_o)
      2'b00: n43916_o = n43911_o;
      2'b01: n43916_o = n43912_o;
      2'b10: n43916_o = n43913_o;
      2'b11: n43916_o = n43914_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n43917_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n43918_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n43919_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n43920_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n43921_o = n42990_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n43921_o)
      2'b00: n43922_o = n43917_o;
      2'b01: n43922_o = n43918_o;
      2'b10: n43922_o = n43919_o;
      2'b11: n43922_o = n43920_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n43923_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n43924_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n43925_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n43926_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n43927_o = n43000_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n43927_o)
      2'b00: n43928_o = n43923_o;
      2'b01: n43928_o = n43924_o;
      2'b10: n43928_o = n43925_o;
      2'b11: n43928_o = n43926_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n43929_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n43930_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n43931_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n43932_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n43933_o = n43010_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n43933_o)
      2'b00: n43934_o = n43929_o;
      2'b01: n43934_o = n43930_o;
      2'b10: n43934_o = n43931_o;
      2'b11: n43934_o = n43932_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n43935_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n43936_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n43937_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n43938_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n43939_o = n43014_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n43939_o)
      2'b00: n43940_o = n43935_o;
      2'b01: n43940_o = n43936_o;
      2'b10: n43940_o = n43937_o;
      2'b11: n43940_o = n43938_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n43941_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n43942_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n43943_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n43944_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n43945_o = n43019_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n43945_o)
      2'b00: n43946_o = n43941_o;
      2'b01: n43946_o = n43942_o;
      2'b10: n43946_o = n43943_o;
      2'b11: n43946_o = n43944_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n43947_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n43948_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n43949_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n43950_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n43951_o = n43027_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n43951_o)
      2'b00: n43952_o = n43947_o;
      2'b01: n43952_o = n43948_o;
      2'b10: n43952_o = n43949_o;
      2'b11: n43952_o = n43950_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n43953_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n43954_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n43955_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n43956_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n43957_o = n43037_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n43957_o)
      2'b00: n43958_o = n43953_o;
      2'b01: n43958_o = n43954_o;
      2'b10: n43958_o = n43955_o;
      2'b11: n43958_o = n43956_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n43959_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n43960_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n43961_o = iregisters_r[38:26];
  assign n43962_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n43963_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n43964_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n43965_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n43966_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n43967_o = n43108_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n43967_o)
      2'b00: n43968_o = n43959_o;
      2'b01: n43968_o = n43960_o;
      2'b10: n43968_o = n43961_o;
      2'b11: n43968_o = n43962_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n43969_o = n43108_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n43969_o)
      2'b00: n43970_o = n43963_o;
      2'b01: n43970_o = n43964_o;
      2'b10: n43970_o = n43965_o;
      2'b11: n43970_o = n43966_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n43971_o = n43108_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n43972_o = n43971_o ? n43970_o : n43968_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n43973_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n43974_o = iregisters_r[25:13];
  assign n43975_o = iregisters_r[38:26];
  assign n43976_o = iregisters_r[51:39];
  assign n43977_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n43978_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n43979_o = iregisters_r[90:78];
  assign n43980_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n43981_o = n43112_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n43981_o)
      2'b00: n43982_o = n43973_o;
      2'b01: n43982_o = n43974_o;
      2'b10: n43982_o = n43975_o;
      2'b11: n43982_o = n43976_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n43983_o = n43112_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n43983_o)
      2'b00: n43984_o = n43977_o;
      2'b01: n43984_o = n43978_o;
      2'b10: n43984_o = n43979_o;
      2'b11: n43984_o = n43980_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n43985_o = n43112_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n43986_o = n43985_o ? n43984_o : n43982_o;
endmodule

module instr_decoder2_1_2
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n41722_o;
  wire n41724_o;
  wire n41727_o;
  wire n41729_o;
  wire n41731_o;
  wire n41733_o;
  wire [5:0] n41734_o;
  wire [3:0] n41736_o;
  wire [3:0] n41738_o;
  wire [3:0] n41739_o;
  wire [3:0] n41740_o;
  reg [3:0] n41741_o;
  wire [8:0] n41743_o;
  wire [8:0] n41745_o;
  wire [8:0] n41746_o;
  wire [8:0] n41747_o;
  reg [8:0] n41748_o;
  wire [12:0] n41751_o;
  wire n41759_o;
  wire n41761_o;
  wire n41764_o;
  wire n41766_o;
  wire n41768_o;
  wire n41770_o;
  wire [5:0] n41771_o;
  wire [3:0] n41773_o;
  wire [3:0] n41775_o;
  wire [3:0] n41776_o;
  wire [3:0] n41777_o;
  reg [3:0] n41778_o;
  wire [8:0] n41780_o;
  wire [8:0] n41782_o;
  wire [8:0] n41783_o;
  wire [8:0] n41784_o;
  reg [8:0] n41785_o;
  wire [12:0] n41788_o;
  wire [7:0] n41789_o;
  wire n41790_o;
  wire [4:0] n41791_o;
  wire [4:0] n41792_o;
  wire [11:0] n41794_o;
  wire [11:0] n41795_o;
  wire [11:0] n41796_o;
  wire [11:0] n41797_o;
  wire [3:0] n41798_o;
  wire [3:0] n41799_o;
  wire [3:0] n41800_o;
  wire [3:0] n41801_o;
  wire n41802_o;
  wire n41803_o;
  wire n41804_o;
  wire n41805_o;
  wire n41808_o;
  wire n41809_o;
  wire n41810_o;
  wire n41811_o;
  wire n41812_o;
  wire n41816_o;
  wire n41817_o;
  wire n41818_o;
  wire n41819_o;
  wire n41820_o;
  wire n41824_o;
  wire n41825_o;
  wire [51:0] n41827_o;
  wire [51:0] n41828_o;
  wire [1:0] n41829_o;
  wire n41833_o;
  wire n41834_o;
  wire n41835_o;
  wire n41836_o;
  wire [12:0] n41837_o;
  wire [1:0] n41839_o;
  wire n41843_o;
  wire n41844_o;
  wire n41845_o;
  wire n41846_o;
  wire [12:0] n41847_o;
  wire [1:0] n41849_o;
  wire n41853_o;
  wire n41854_o;
  wire n41855_o;
  wire n41856_o;
  wire [12:0] n41857_o;
  wire [1:0] n41859_o;
  wire [1:0] n41863_o;
  wire [1:0] n41868_o;
  wire [1:0] n41876_o;
  wire n41880_o;
  wire n41881_o;
  wire n41882_o;
  wire n41883_o;
  wire [12:0] n41884_o;
  wire [1:0] n41886_o;
  wire n41890_o;
  wire n41891_o;
  wire [12:0] n41892_o;
  wire n41893_o;
  wire [7:0] n41894_o;
  wire [7:0] n41895_o;
  wire n41898_o;
  wire [51:0] n41900_o;
  wire [25:0] n41901_o;
  wire n41902_o;
  wire n41903_o;
  wire [12:0] n41904_o;
  wire [12:0] n41905_o;
  wire [12:0] n41906_o;
  wire n41907_o;
  wire n41908_o;
  wire [12:0] n41909_o;
  wire [12:0] n41910_o;
  wire [12:0] n41911_o;
  wire [103:0] n41922_o;
  wire [4:0] n41947_o;
  wire [3:0] n41948_o;
  wire [3:0] n41949_o;
  wire [3:0] n41950_o;
  wire [12:0] n41951_o;
  wire n41955_o;
  wire [2:0] n41957_o;
  wire [2:0] n41961_o;
  wire n41966_o;
  wire n41967_o;
  wire n41969_o;
  wire [2:0] n41970_o;
  wire [2:0] n41972_o;
  wire n41975_o;
  wire n41977_o;
  wire n41980_o;
  wire n41982_o;
  wire [2:0] n41984_o;
  wire n41986_o;
  wire n41988_o;
  wire [2:0] n41990_o;
  wire n41992_o;
  wire [4:0] n41994_o;
  wire [1:0] n42142_o;
  wire n42144_o;
  wire n42146_o;
  wire n42147_o;
  wire [2:0] n42148_o;
  wire [12:0] n42160_o;
  wire [12:0] n42161_o;
  wire [12:0] n42162_o;
  wire [9:0] n42164_o;
  wire [12:0] n42168_o;
  wire [12:0] n42169_o;
  wire [12:0] n42171_o;
  wire [9:0] n42173_o;
  wire [12:0] n42177_o;
  wire [12:0] n42178_o;
  wire n42180_o;
  wire [1:0] n42181_o;
  wire n42183_o;
  wire n42184_o;
  wire [11:0] n42185_o;
  wire [8:0] n42186_o;
  wire [8:0] n42187_o;
  wire [2:0] n42188_o;
  wire [2:0] n42189_o;
  wire [2:0] n42190_o;
  wire n42192_o;
  wire [1:0] n42193_o;
  wire n42195_o;
  wire n42196_o;
  wire n42198_o;
  wire n42199_o;
  wire n42201_o;
  wire [4:0] n42202_o;
  wire [8:0] n42203_o;
  wire [4:0] n42204_o;
  wire [5:0] n42206_o;
  wire [2:0] n42207_o;
  wire [8:0] n42208_o;
  wire [8:0] n42209_o;
  wire [2:0] n42210_o;
  wire [12:0] n42211_o;
  wire n42212_o;
  wire [11:0] n42213_o;
  wire [8:0] n42214_o;
  wire [8:0] n42215_o;
  wire [2:0] n42216_o;
  wire n42218_o;
  wire [4:0] n42219_o;
  wire [8:0] n42220_o;
  wire [4:0] n42221_o;
  wire [5:0] n42223_o;
  wire [2:0] n42224_o;
  wire [8:0] n42225_o;
  wire [8:0] n42226_o;
  wire [2:0] n42227_o;
  wire [11:0] n42228_o;
  wire [11:0] n42229_o;
  wire [11:0] n42230_o;
  wire [11:0] n42231_o;
  wire [11:0] n42232_o;
  wire [11:0] n42235_o;
  wire [11:0] n42236_o;
  wire [1:0] n42252_o;
  wire n42254_o;
  wire n42256_o;
  wire n42257_o;
  wire [2:0] n42258_o;
  wire [12:0] n42270_o;
  wire [12:0] n42271_o;
  wire [12:0] n42272_o;
  wire [9:0] n42274_o;
  wire [12:0] n42278_o;
  wire [12:0] n42279_o;
  wire [12:0] n42281_o;
  wire [9:0] n42283_o;
  wire [12:0] n42287_o;
  wire [12:0] n42288_o;
  wire n42290_o;
  wire [1:0] n42291_o;
  wire n42293_o;
  wire n42294_o;
  wire [11:0] n42295_o;
  wire [8:0] n42296_o;
  wire [8:0] n42297_o;
  wire [2:0] n42298_o;
  wire [2:0] n42299_o;
  wire [2:0] n42300_o;
  wire n42302_o;
  wire [1:0] n42303_o;
  wire n42305_o;
  wire n42306_o;
  wire n42308_o;
  wire n42309_o;
  wire n42311_o;
  wire [4:0] n42312_o;
  wire [8:0] n42313_o;
  wire [4:0] n42314_o;
  wire [5:0] n42316_o;
  wire [2:0] n42317_o;
  wire [8:0] n42318_o;
  wire [8:0] n42319_o;
  wire [2:0] n42320_o;
  wire [12:0] n42321_o;
  wire n42322_o;
  wire [11:0] n42323_o;
  wire [8:0] n42324_o;
  wire [8:0] n42325_o;
  wire [2:0] n42326_o;
  wire n42328_o;
  wire [4:0] n42329_o;
  wire [8:0] n42330_o;
  wire [4:0] n42331_o;
  wire [5:0] n42333_o;
  wire [2:0] n42334_o;
  wire [8:0] n42335_o;
  wire [8:0] n42336_o;
  wire [2:0] n42337_o;
  wire [11:0] n42338_o;
  wire [11:0] n42339_o;
  wire [11:0] n42340_o;
  wire [11:0] n42341_o;
  wire [11:0] n42342_o;
  wire [11:0] n42345_o;
  wire [11:0] n42346_o;
  wire [1:0] n42362_o;
  wire n42364_o;
  wire n42366_o;
  wire n42367_o;
  wire [2:0] n42368_o;
  wire [12:0] n42380_o;
  wire [12:0] n42381_o;
  wire [12:0] n42382_o;
  wire [9:0] n42384_o;
  wire [12:0] n42388_o;
  wire [12:0] n42389_o;
  wire [12:0] n42391_o;
  wire [9:0] n42393_o;
  wire [12:0] n42397_o;
  wire [12:0] n42398_o;
  wire n42400_o;
  wire [1:0] n42401_o;
  wire n42403_o;
  wire n42404_o;
  wire [11:0] n42405_o;
  wire [8:0] n42406_o;
  wire [8:0] n42407_o;
  wire [2:0] n42408_o;
  wire [2:0] n42409_o;
  wire [2:0] n42410_o;
  wire n42412_o;
  wire [1:0] n42413_o;
  wire n42415_o;
  wire n42416_o;
  wire n42418_o;
  wire n42419_o;
  wire n42421_o;
  wire [4:0] n42422_o;
  wire [8:0] n42423_o;
  wire [4:0] n42424_o;
  wire [5:0] n42426_o;
  wire [2:0] n42427_o;
  wire [8:0] n42428_o;
  wire [8:0] n42429_o;
  wire [2:0] n42430_o;
  wire [12:0] n42431_o;
  wire n42432_o;
  wire [11:0] n42433_o;
  wire [8:0] n42434_o;
  wire [8:0] n42435_o;
  wire [2:0] n42436_o;
  wire n42438_o;
  wire [4:0] n42439_o;
  wire [8:0] n42440_o;
  wire [4:0] n42441_o;
  wire [5:0] n42443_o;
  wire [2:0] n42444_o;
  wire [8:0] n42445_o;
  wire [8:0] n42446_o;
  wire [2:0] n42447_o;
  wire [11:0] n42448_o;
  wire [11:0] n42449_o;
  wire [11:0] n42450_o;
  wire [11:0] n42451_o;
  wire [11:0] n42452_o;
  wire [11:0] n42455_o;
  wire [11:0] n42456_o;
  wire [1:0] n42472_o;
  wire n42474_o;
  wire n42476_o;
  wire n42477_o;
  wire [2:0] n42478_o;
  wire [12:0] n42490_o;
  wire [12:0] n42491_o;
  wire [12:0] n42492_o;
  wire [9:0] n42494_o;
  wire [12:0] n42498_o;
  wire [12:0] n42499_o;
  wire [12:0] n42501_o;
  wire [9:0] n42503_o;
  wire [12:0] n42507_o;
  wire [12:0] n42508_o;
  wire n42510_o;
  wire [1:0] n42511_o;
  wire n42513_o;
  wire n42514_o;
  wire [11:0] n42515_o;
  wire [8:0] n42516_o;
  wire [8:0] n42517_o;
  wire [2:0] n42518_o;
  wire [2:0] n42519_o;
  wire [2:0] n42520_o;
  wire n42522_o;
  wire [1:0] n42523_o;
  wire n42525_o;
  wire n42526_o;
  wire n42528_o;
  wire n42529_o;
  wire n42531_o;
  wire [4:0] n42532_o;
  wire [8:0] n42533_o;
  wire [4:0] n42534_o;
  wire [5:0] n42536_o;
  wire [2:0] n42537_o;
  wire [8:0] n42538_o;
  wire [8:0] n42539_o;
  wire [2:0] n42540_o;
  wire [12:0] n42541_o;
  wire n42542_o;
  wire [11:0] n42543_o;
  wire [8:0] n42544_o;
  wire [8:0] n42545_o;
  wire [2:0] n42546_o;
  wire n42548_o;
  wire [4:0] n42549_o;
  wire [8:0] n42550_o;
  wire [4:0] n42551_o;
  wire [5:0] n42553_o;
  wire [2:0] n42554_o;
  wire [8:0] n42555_o;
  wire [8:0] n42556_o;
  wire [2:0] n42557_o;
  wire [11:0] n42558_o;
  wire [11:0] n42559_o;
  wire [11:0] n42560_o;
  wire [11:0] n42561_o;
  wire [11:0] n42562_o;
  wire [11:0] n42565_o;
  wire [11:0] n42566_o;
  wire n42573_o;
  wire [11:0] n42575_o;
  wire [6:0] n42576_o;
  wire [7:0] n42577_o;
  wire [3:0] n42579_o;
  wire [7:0] n42580_o;
  wire [6:0] n42581_o;
  wire [7:0] n42582_o;
  wire [7:0] n42583_o;
  wire n42586_o;
  wire n42588_o;
  wire n42590_o;
  wire n42592_o;
  wire n42594_o;
  wire [4:0] n42596_o;
  wire [7:0] n42601_o;
  wire [7:0] n42603_o;
  wire [7:0] n42605_o;
  wire [7:0] n42607_o;
  reg [3:0] n42678_q;
  reg [3:0] n42679_q;
  reg [3:0] n42680_q;
  reg [3:0] n42681_q;
  reg [3:0] n42682_q;
  reg [3:0] n42683_q;
  reg n42685_q;
  reg n42686_q;
  reg [12:0] n42687_q;
  reg [12:0] n42688_q;
  reg [12:0] n42689_q;
  reg n42690_q;
  reg n42691_q;
  reg n42692_q;
  reg n42693_q;
  reg n42695_q;
  reg n42696_q;
  reg n42697_q;
  reg n42698_q;
  reg n42699_q;
  reg n42700_q;
  reg [11:0] n42701_q;
  reg n42702_q;
  reg n42703_q;
  reg n42704_q;
  reg [4:0] n42705_q;
  wire [11:0] n42706_o;
  reg [11:0] n42707_q;
  wire [11:0] n42708_o;
  reg [11:0] n42709_q;
  wire [11:0] n42710_o;
  reg [11:0] n42711_q;
  reg n42712_q;
  reg n42713_q;
  reg n42714_q;
  reg n42715_q;
  reg n42716_q;
  reg n42717_q;
  reg [4:0] n42719_q;
  reg [3:0] n42720_q;
  reg [3:0] n42721_q;
  reg [3:0] n42722_q;
  reg [12:0] n42723_q;
  reg [4:0] n42724_q;
  reg [3:0] n42725_q;
  reg [3:0] n42726_q;
  reg [3:0] n42727_q;
  reg [3:0] n42728_q;
  reg [3:0] n42729_q;
  reg [12:0] n42730_q;
  reg [12:0] n42731_q;
  reg [2:0] n42732_q;
  reg [2:0] n42733_q;
  reg [2:0] n42734_q;
  reg [2:0] n42735_q;
  reg n42737_q;
  reg n42738_q;
  reg n42739_q;
  reg n42740_q;
  reg [4:0] n42742_q;
  reg [103:0] n42743_q;
  reg [12:0] n42744_q;
  reg [12:0] n42745_q;
  reg [12:0] n42746_q;
  reg [12:0] n42747_q;
  reg [12:0] n42748_q;
  reg [12:0] n42749_q;
  reg [7:0] n42750_q;
  reg [7:0] n42751_q;
  reg [7:0] n42752_q;
  reg [7:0] n42753_q;
  reg [7:0] n42754_q;
  reg [7:0] n42755_q;
  reg [7:0] n42756_q;
  reg [7:0] n42757_q;
  reg [7:0] n42758_q;
  reg [12:0] n42759_q;
  wire [12:0] n42760_o;
  wire [12:0] n42761_o;
  wire [12:0] n42762_o;
  wire [12:0] n42763_o;
  wire [1:0] n42764_o;
  reg [12:0] n42765_o;
  wire [12:0] n42766_o;
  wire [12:0] n42767_o;
  wire [12:0] n42768_o;
  wire [12:0] n42769_o;
  wire [1:0] n42770_o;
  reg [12:0] n42771_o;
  wire [12:0] n42772_o;
  wire [12:0] n42773_o;
  wire [12:0] n42774_o;
  wire [12:0] n42775_o;
  wire [1:0] n42776_o;
  reg [12:0] n42777_o;
  wire [12:0] n42778_o;
  wire [12:0] n42779_o;
  wire [12:0] n42780_o;
  wire [12:0] n42781_o;
  wire [1:0] n42782_o;
  reg [12:0] n42783_o;
  wire [12:0] n42784_o;
  wire [12:0] n42785_o;
  wire [12:0] n42786_o;
  wire [12:0] n42787_o;
  wire [1:0] n42788_o;
  reg [12:0] n42789_o;
  wire [12:0] n42790_o;
  wire [12:0] n42791_o;
  wire [12:0] n42792_o;
  wire [12:0] n42793_o;
  wire [1:0] n42794_o;
  reg [12:0] n42795_o;
  wire [12:0] n42796_o;
  wire [12:0] n42797_o;
  wire [12:0] n42798_o;
  wire [12:0] n42799_o;
  wire [1:0] n42800_o;
  reg [12:0] n42801_o;
  wire [12:0] n42802_o;
  wire [12:0] n42803_o;
  wire [12:0] n42804_o;
  wire [12:0] n42805_o;
  wire [1:0] n42806_o;
  reg [12:0] n42807_o;
  wire [12:0] n42808_o;
  wire [12:0] n42809_o;
  wire [12:0] n42810_o;
  wire [12:0] n42811_o;
  wire [12:0] n42812_o;
  wire [12:0] n42813_o;
  wire [12:0] n42814_o;
  wire [12:0] n42815_o;
  wire [1:0] n42816_o;
  reg [12:0] n42817_o;
  wire [1:0] n42818_o;
  reg [12:0] n42819_o;
  wire n42820_o;
  wire [12:0] n42821_o;
  wire [12:0] n42822_o;
  wire [12:0] n42823_o;
  wire [12:0] n42824_o;
  wire [12:0] n42825_o;
  wire [12:0] n42826_o;
  wire [12:0] n42827_o;
  wire [12:0] n42828_o;
  wire [12:0] n42829_o;
  wire [1:0] n42830_o;
  reg [12:0] n42831_o;
  wire [1:0] n42832_o;
  reg [12:0] n42833_o;
  wire n42834_o;
  wire [12:0] n42835_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n41894_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n41751_o;
  assign i_x2_out = n41788_o;
  assign result_waddr_out = n41789_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n42678_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n42679_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n42680_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n42681_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n42682_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n42683_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n42685_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n42686_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n42687_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n42688_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n42689_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n42690_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n42691_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n42692_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n42693_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n41792_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n42695_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n42696_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n41790_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n42697_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n41812_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n42698_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n41820_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n42699_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n41825_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n42700_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n42701_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n41794_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n41795_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n41796_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n41797_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n41798_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n41799_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n41800_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n41801_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n41802_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n41803_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n41804_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n41805_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n42702_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n42703_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n42704_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n42705_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n42707_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n42709_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n42711_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n42236_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n42346_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n42456_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n42566_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n42712_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n42713_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n42714_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n42715_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n42716_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n42717_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n41947_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n41948_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n41949_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n41950_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n41951_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n42719_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n42720_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n42721_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n42722_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n42723_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n42724_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n42725_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n42726_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n42727_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n42728_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n42729_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n42730_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n42731_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n42732_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n42733_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n42734_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n42735_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n42737_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n42738_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n42739_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n42740_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n42742_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n42743_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n41827_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n41828_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n42744_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n42745_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n42746_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n42747_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n42748_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n42749_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n41837_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n41847_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n41857_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n42783_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n42789_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n42795_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n41892_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n41884_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n42807_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n42750_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n42751_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n42752_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n42753_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n42754_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n42755_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n42756_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n42757_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n42758_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n42759_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n41722_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n41724_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n41727_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n41729_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n41731_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n41733_o = imu_x1_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41734_o = {n41733_o, n41731_o, n41729_o, n41727_o, n41724_o, n41722_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41736_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41738_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41739_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41740_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n41734_o)
      6'b100000: n41741_o = n41739_o;
      6'b010000: n41741_o = n41738_o;
      6'b001000: n41741_o = 4'b0110;
      6'b000100: n41741_o = instruction_tid_rrr;
      6'b000010: n41741_o = n41736_o;
      6'b000001: n41741_o = 4'b0000;
      default: n41741_o = n41740_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41743_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41745_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41746_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41747_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n41734_o)
      6'b100000: n41748_o = n41746_o;
      6'b010000: n41748_o = n41745_o;
      6'b001000: n41748_o = 9'b000000000;
      6'b000100: n41748_o = 9'b000000000;
      6'b000010: n41748_o = n41743_o;
      6'b000001: n41748_o = 9'b000000000;
      default: n41748_o = n41747_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41751_o = {n41748_o, n41741_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n41759_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n41761_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n41764_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n41766_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n41768_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n41770_o = imu_x2_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41771_o = {n41770_o, n41768_o, n41766_o, n41764_o, n41761_o, n41759_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41773_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41775_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41776_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n41777_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n41771_o)
      6'b100000: n41778_o = n41776_o;
      6'b010000: n41778_o = n41775_o;
      6'b001000: n41778_o = 4'b0110;
      6'b000100: n41778_o = instruction_tid_rrr;
      6'b000010: n41778_o = n41773_o;
      6'b000001: n41778_o = 4'b0000;
      default: n41778_o = n41777_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41780_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41782_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41783_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41784_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n41771_o)
      6'b100000: n41785_o = n41783_o;
      6'b010000: n41785_o = n41782_o;
      6'b001000: n41785_o = 9'b000000000;
      6'b000100: n41785_o = 9'b000000000;
      6'b000010: n41785_o = n41780_o;
      6'b000001: n41785_o = 9'b000000000;
      default: n41785_o = n41784_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n41788_o = {n41785_o, n41778_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n41789_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n41790_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n41791_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n41792_o = instruction_mu_valid_in ? n41791_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n41794_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n41795_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n41796_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n41797_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n41798_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n41799_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n41800_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n41801_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n41802_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n41803_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n41804_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n41805_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n41808_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n41809_o = n41808_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n41810_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n41811_o = n41810_o & n41809_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n41812_o = n41811_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n41816_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n41817_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n41818_o = n41817_o & n41816_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n41819_o = n41818_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n41820_o = n41819_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n41824_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n41825_o = n41824_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n41827_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n41828_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n41829_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n41833_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n41834_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n41835_o = ~n41834_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n41836_o = n41833_o | n41835_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n41837_o = n41836_o ? n42765_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n41839_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n41843_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n41844_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n41845_o = ~n41844_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n41846_o = n41843_o | n41845_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n41847_o = n41846_o ? n42771_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n41849_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n41853_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n41854_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n41855_o = ~n41854_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n41856_o = n41853_o | n41855_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n41857_o = n41856_o ? n42777_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n41859_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n41863_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n41868_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n41876_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n41880_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n41881_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n41882_o = ~n41881_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n41883_o = n41880_o | n41882_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n41884_o = n41883_o ? n42801_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n41886_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n41890_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n41891_o = ~n41890_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n41892_o = n41891_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n41893_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n41894_o = n41893_o ? mu_lane_rrrrrr : n41895_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n41895_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n41898_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n41900_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n41901_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n41902_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n41903_o = ~n41902_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n41904_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n41905_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n41906_o = n41903_o ? n41904_o : n41905_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n41907_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n41908_o = ~n41907_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n41909_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n41910_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n41911_o = n41908_o ? n41909_o : n41910_o;
  assign n41922_o = {n41900_o, n41906_o, n41911_o, n41901_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n41947_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n41948_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n41949_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n41950_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n41951_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n41955_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n41957_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n41961_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n41966_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n41967_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n41969_o = n41967_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n41970_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n41972_o = n41969_o ? n41970_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n41975_o = n41969_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n41977_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n41980_o = n41977_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n41982_o = n41966_o ? n41980_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n41984_o = n41966_o ? n41972_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n41986_o = n41966_o ? n41975_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n41988_o = got_imu_rr ? n41982_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n41990_o = got_imu_rr ? n41984_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n41992_o = got_imu_rr ? n41986_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n41994_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n42142_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n42144_o = n42142_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n42146_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n42147_o = n42144_o | n42146_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n42148_o = mu_x1_parm1[2:0];
  assign n42160_o = {1'b0, mu_x1_parm1};
  assign n42161_o = {10'b0000000000, n42148_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n42162_o = n42147_o ? n42161_o : n42160_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n42164_o = mu_x1_i1_1[9:0];
  assign n42168_o = {n42164_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n42169_o = mu_x1_vector ? n42168_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n42171_o = mu_x1_i0_1 + n42162_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n42173_o = n42171_o[9:0];
  assign n42177_o = {n42173_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42178_o = mu_x1_vector ? n42177_o : n42171_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n42180_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n42181_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n42183_o = n42181_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n42184_o = n42180_o | n42183_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n42185_o = n42178_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n42186_o = n42185_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n42187_o = ~n42186_o;
  assign n42188_o = n42177_o[2:0];
  assign n42189_o = n42171_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42190_o = mu_x1_vector ? n42188_o : n42189_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n42192_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n42193_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n42195_o = n42193_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n42196_o = n42192_o | n42195_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n42198_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n42199_o = n42196_o | n42198_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n42201_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n42202_o = n42178_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n42203_o = {n42202_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n42204_o = n42178_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n42206_o = {1'b0, n42204_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n42207_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n42208_o = {n42206_o, n42207_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n42209_o = n42201_o ? n42203_o : n42208_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n42210_o = n42178_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n42211_o = n42169_o + n42178_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n42212_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n42213_o = n42211_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n42214_o = n42213_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n42215_o = ~n42214_o;
  assign n42216_o = n42211_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n42218_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n42219_o = n42211_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n42220_o = {n42219_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n42221_o = n42211_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n42223_o = {1'b0, n42221_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n42224_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n42225_o = {n42223_o, n42224_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n42226_o = n42218_o ? n42220_o : n42225_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n42227_o = n42211_o[2:0];
  assign n42228_o = {n42226_o, n42227_o};
  assign n42229_o = {n42215_o, n42216_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n42230_o = n42212_o ? n42229_o : n42228_o;
  assign n42231_o = {n42209_o, n42210_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n42232_o = n42199_o ? n42231_o : n42230_o;
  assign n42235_o = {n42187_o, n42190_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n42236_o = n42184_o ? n42235_o : n42232_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n42252_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n42254_o = n42252_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n42256_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n42257_o = n42254_o | n42256_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n42258_o = mu_x2_parm1[2:0];
  assign n42270_o = {1'b0, mu_x2_parm1};
  assign n42271_o = {10'b0000000000, n42258_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n42272_o = n42257_o ? n42271_o : n42270_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n42274_o = mu_x2_i1_1[9:0];
  assign n42278_o = {n42274_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n42279_o = mu_x2_vector ? n42278_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n42281_o = mu_x2_i0_1 + n42272_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n42283_o = n42281_o[9:0];
  assign n42287_o = {n42283_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42288_o = mu_x2_vector ? n42287_o : n42281_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n42290_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n42291_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n42293_o = n42291_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n42294_o = n42290_o | n42293_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n42295_o = n42288_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n42296_o = n42295_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n42297_o = ~n42296_o;
  assign n42298_o = n42287_o[2:0];
  assign n42299_o = n42281_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42300_o = mu_x2_vector ? n42298_o : n42299_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n42302_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n42303_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n42305_o = n42303_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n42306_o = n42302_o | n42305_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n42308_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n42309_o = n42306_o | n42308_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n42311_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n42312_o = n42288_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n42313_o = {n42312_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n42314_o = n42288_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n42316_o = {1'b0, n42314_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n42317_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n42318_o = {n42316_o, n42317_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n42319_o = n42311_o ? n42313_o : n42318_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n42320_o = n42288_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n42321_o = n42279_o + n42288_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n42322_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n42323_o = n42321_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n42324_o = n42323_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n42325_o = ~n42324_o;
  assign n42326_o = n42321_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n42328_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n42329_o = n42321_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n42330_o = {n42329_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n42331_o = n42321_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n42333_o = {1'b0, n42331_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n42334_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n42335_o = {n42333_o, n42334_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n42336_o = n42328_o ? n42330_o : n42335_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n42337_o = n42321_o[2:0];
  assign n42338_o = {n42336_o, n42337_o};
  assign n42339_o = {n42325_o, n42326_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n42340_o = n42322_o ? n42339_o : n42338_o;
  assign n42341_o = {n42319_o, n42320_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n42342_o = n42309_o ? n42341_o : n42340_o;
  assign n42345_o = {n42297_o, n42300_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n42346_o = n42294_o ? n42345_o : n42342_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n42362_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n42364_o = n42362_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n42366_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n42367_o = n42364_o | n42366_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n42368_o = mu_x3_parm1[2:0];
  assign n42380_o = {1'b0, mu_x3_parm1};
  assign n42381_o = {10'b0000000000, n42368_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n42382_o = n42367_o ? n42381_o : n42380_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n42384_o = mu_x3_i1_1[9:0];
  assign n42388_o = {n42384_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n42389_o = mu_x3_vector ? n42388_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n42391_o = mu_x3_i0_1 + n42382_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n42393_o = n42391_o[9:0];
  assign n42397_o = {n42393_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42398_o = mu_x3_vector ? n42397_o : n42391_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n42400_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n42401_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n42403_o = n42401_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n42404_o = n42400_o | n42403_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n42405_o = n42398_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n42406_o = n42405_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n42407_o = ~n42406_o;
  assign n42408_o = n42397_o[2:0];
  assign n42409_o = n42391_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42410_o = mu_x3_vector ? n42408_o : n42409_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n42412_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n42413_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n42415_o = n42413_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n42416_o = n42412_o | n42415_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n42418_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n42419_o = n42416_o | n42418_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n42421_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n42422_o = n42398_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n42423_o = {n42422_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n42424_o = n42398_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n42426_o = {1'b0, n42424_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n42427_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n42428_o = {n42426_o, n42427_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n42429_o = n42421_o ? n42423_o : n42428_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n42430_o = n42398_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n42431_o = n42389_o + n42398_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n42432_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n42433_o = n42431_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n42434_o = n42433_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n42435_o = ~n42434_o;
  assign n42436_o = n42431_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n42438_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n42439_o = n42431_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n42440_o = {n42439_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n42441_o = n42431_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n42443_o = {1'b0, n42441_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n42444_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n42445_o = {n42443_o, n42444_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n42446_o = n42438_o ? n42440_o : n42445_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n42447_o = n42431_o[2:0];
  assign n42448_o = {n42446_o, n42447_o};
  assign n42449_o = {n42435_o, n42436_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n42450_o = n42432_o ? n42449_o : n42448_o;
  assign n42451_o = {n42429_o, n42430_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n42452_o = n42419_o ? n42451_o : n42450_o;
  assign n42455_o = {n42407_o, n42410_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n42456_o = n42404_o ? n42455_o : n42452_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n42472_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n42474_o = n42472_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n42476_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n42477_o = n42474_o | n42476_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n42478_o = mu_y_parm1[2:0];
  assign n42490_o = {1'b0, mu_y_parm1};
  assign n42491_o = {10'b0000000000, n42478_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n42492_o = n42477_o ? n42491_o : n42490_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n42494_o = mu_y_i1_1[9:0];
  assign n42498_o = {n42494_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n42499_o = mu_y_vector ? n42498_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n42501_o = mu_y_i0_1 + n42492_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n42503_o = n42501_o[9:0];
  assign n42507_o = {n42503_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42508_o = mu_y_vector ? n42507_o : n42501_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n42510_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n42511_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n42513_o = n42511_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n42514_o = n42510_o | n42513_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n42515_o = n42508_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n42516_o = n42515_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n42517_o = ~n42516_o;
  assign n42518_o = n42507_o[2:0];
  assign n42519_o = n42501_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n42520_o = mu_y_vector ? n42518_o : n42519_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n42522_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n42523_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n42525_o = n42523_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n42526_o = n42522_o | n42525_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n42528_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n42529_o = n42526_o | n42528_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n42531_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n42532_o = n42508_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n42533_o = {n42532_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n42534_o = n42508_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n42536_o = {1'b0, n42534_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n42537_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n42538_o = {n42536_o, n42537_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n42539_o = n42531_o ? n42533_o : n42538_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n42540_o = n42508_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n42541_o = n42499_o + n42508_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n42542_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n42543_o = n42541_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n42544_o = n42543_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n42545_o = ~n42544_o;
  assign n42546_o = n42541_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n42548_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n42549_o = n42541_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n42550_o = {n42549_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n42551_o = n42541_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n42553_o = {1'b0, n42551_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n42554_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n42555_o = {n42553_o, n42554_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n42556_o = n42548_o ? n42550_o : n42555_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n42557_o = n42541_o[2:0];
  assign n42558_o = {n42556_o, n42557_o};
  assign n42559_o = {n42545_o, n42546_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n42560_o = n42542_o ? n42559_o : n42558_o;
  assign n42561_o = {n42539_o, n42540_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n42562_o = n42529_o ? n42561_o : n42560_o;
  assign n42565_o = {n42517_o, n42520_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n42566_o = n42514_o ? n42565_o : n42562_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n42573_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n42575_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n42576_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n42577_o = {instruction_vm_in, n42576_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n42579_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n42580_o = {n42579_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n42581_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n42582_o = {instruction_vm_in, n42581_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n42583_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42586_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42588_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42590_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42592_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42594_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42596_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42601_o = instruction_tid_valid_in ? n42583_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42603_o = instruction_tid_valid_in ? n42582_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42605_o = instruction_tid_valid_in ? n42580_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n42607_o = instruction_tid_valid_in ? n42577_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42678_q <= 4'b0000;
    else
      n42678_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42679_q <= 4'b0000;
    else
      n42679_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42680_q <= 4'b0000;
    else
      n42680_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42681_q <= 4'b0000;
    else
      n42681_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42682_q <= 4'b0000;
    else
      n42682_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42683_q <= 4'b0000;
    else
      n42683_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42685_q <= 1'b0;
    else
      n42685_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42686_q <= 1'b0;
    else
      n42686_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42687_q <= 13'b0000000000000;
    else
      n42687_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42688_q <= 13'b0000000000000;
    else
      n42688_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42689_q <= 13'b0000000000000;
    else
      n42689_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42690_q <= 1'b0;
    else
      n42690_q <= n41988_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42691_q <= 1'b0;
    else
      n42691_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42692_q <= 1'b0;
    else
      n42692_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42693_q <= 1'b0;
    else
      n42693_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42695_q <= 1'b0;
    else
      n42695_q <= n42586_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42696_q <= 1'b0;
    else
      n42696_q <= n42588_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42697_q <= 1'b0;
    else
      n42697_q <= n42590_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42698_q <= 1'b0;
    else
      n42698_q <= n42592_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42699_q <= 1'b0;
    else
      n42699_q <= n42594_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42700_q <= 1'b0;
    else
      n42700_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42701_q <= 12'b000000000000;
    else
      n42701_q <= n42575_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42702_q <= 1'b0;
    else
      n42702_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42703_q <= 1'b0;
    else
      n42703_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42704_q <= 1'b0;
    else
      n42704_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42705_q <= 5'b00000;
    else
      n42705_q <= n42596_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n42706_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42707_q <= 12'b000000000000;
    else
      n42707_q <= n42706_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n42708_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42709_q <= 12'b000000000000;
    else
      n42709_q <= n42708_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n42710_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42711_q <= 12'b000000000000;
    else
      n42711_q <= n42710_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42712_q <= 1'b0;
    else
      n42712_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42713_q <= 1'b0;
    else
      n42713_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42714_q <= 1'b0;
    else
      n42714_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42715_q <= 1'b0;
    else
      n42715_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42716_q <= 1'b0;
    else
      n42716_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42717_q <= 1'b0;
    else
      n42717_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42719_q <= 5'b00000;
    else
      n42719_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42720_q <= 4'b0000;
    else
      n42720_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42721_q <= 4'b0000;
    else
      n42721_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42722_q <= 4'b0000;
    else
      n42722_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42723_q <= 13'b0000000000000;
    else
      n42723_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42724_q <= 5'b00000;
    else
      n42724_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42725_q <= 4'b0000;
    else
      n42725_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42726_q <= 4'b0000;
    else
      n42726_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42727_q <= 4'b0000;
    else
      n42727_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42728_q <= 4'b0000;
    else
      n42728_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42729_q <= 4'b0000;
    else
      n42729_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42730_q <= 13'b0000000000000;
    else
      n42730_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42731_q <= 13'b0000000000000;
    else
      n42731_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42732_q <= 3'b000;
    else
      n42732_q <= n41990_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42733_q <= 3'b000;
    else
      n42733_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42734_q <= 3'b000;
    else
      n42734_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42735_q <= 3'b000;
    else
      n42735_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42737_q <= 1'b0;
    else
      n42737_q <= n41992_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42738_q <= 1'b0;
    else
      n42738_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42739_q <= 1'b0;
    else
      n42739_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42740_q <= 1'b0;
    else
      n42740_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42742_q <= 5'b00000;
    else
      n42742_q <= n41994_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n41898_o)
    if (n41898_o)
      n42743_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n42743_q <= n41922_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42744_q <= 13'b0000000000000;
    else
      n42744_q <= n42821_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42745_q <= 13'b0000000000000;
    else
      n42745_q <= n42835_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42746_q <= 13'b0000000000000;
    else
      n42746_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42747_q <= 13'b0000000000000;
    else
      n42747_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42748_q <= 13'b0000000000000;
    else
      n42748_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42749_q <= 13'b0000000000000;
    else
      n42749_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42750_q <= 8'b00000000;
    else
      n42750_q <= n42601_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42751_q <= 8'b00000000;
    else
      n42751_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42752_q <= 8'b00000000;
    else
      n42752_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42753_q <= 8'b00000000;
    else
      n42753_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42754_q <= 8'b00000000;
    else
      n42754_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42755_q <= 8'b00000000;
    else
      n42755_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42756_q <= 8'b00000000;
    else
      n42756_q <= n42603_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42757_q <= 8'b00000000;
    else
      n42757_q <= n42605_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n42573_o)
    if (n42573_o)
      n42758_q <= 8'b00000000;
    else
      n42758_q <= n42607_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n41955_o)
    if (n41955_o)
      n42759_q <= 13'b0000000000000;
    else
      n42759_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n42760_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n42761_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n42762_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n42763_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n42764_o = n41829_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n42764_o)
      2'b00: n42765_o = n42760_o;
      2'b01: n42765_o = n42761_o;
      2'b10: n42765_o = n42762_o;
      2'b11: n42765_o = n42763_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n42766_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n42767_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n42768_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n42769_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n42770_o = n41839_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n42770_o)
      2'b00: n42771_o = n42766_o;
      2'b01: n42771_o = n42767_o;
      2'b10: n42771_o = n42768_o;
      2'b11: n42771_o = n42769_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n42772_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n42773_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n42774_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n42775_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n42776_o = n41849_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n42776_o)
      2'b00: n42777_o = n42772_o;
      2'b01: n42777_o = n42773_o;
      2'b10: n42777_o = n42774_o;
      2'b11: n42777_o = n42775_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n42778_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n42779_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n42780_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n42781_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n42782_o = n41859_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n42782_o)
      2'b00: n42783_o = n42778_o;
      2'b01: n42783_o = n42779_o;
      2'b10: n42783_o = n42780_o;
      2'b11: n42783_o = n42781_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n42784_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n42785_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n42786_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n42787_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n42788_o = n41863_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n42788_o)
      2'b00: n42789_o = n42784_o;
      2'b01: n42789_o = n42785_o;
      2'b10: n42789_o = n42786_o;
      2'b11: n42789_o = n42787_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n42790_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n42791_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n42792_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n42793_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n42794_o = n41868_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n42794_o)
      2'b00: n42795_o = n42790_o;
      2'b01: n42795_o = n42791_o;
      2'b10: n42795_o = n42792_o;
      2'b11: n42795_o = n42793_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n42796_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n42797_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n42798_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n42799_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n42800_o = n41876_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n42800_o)
      2'b00: n42801_o = n42796_o;
      2'b01: n42801_o = n42797_o;
      2'b10: n42801_o = n42798_o;
      2'b11: n42801_o = n42799_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n42802_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n42803_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n42804_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n42805_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n42806_o = n41886_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n42806_o)
      2'b00: n42807_o = n42802_o;
      2'b01: n42807_o = n42803_o;
      2'b10: n42807_o = n42804_o;
      2'b11: n42807_o = n42805_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n42808_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n42809_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n42810_o = iregisters_r[38:26];
  assign n42811_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n42812_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n42813_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n42814_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n42815_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n42816_o = n41957_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n42816_o)
      2'b00: n42817_o = n42808_o;
      2'b01: n42817_o = n42809_o;
      2'b10: n42817_o = n42810_o;
      2'b11: n42817_o = n42811_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n42818_o = n41957_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n42818_o)
      2'b00: n42819_o = n42812_o;
      2'b01: n42819_o = n42813_o;
      2'b10: n42819_o = n42814_o;
      2'b11: n42819_o = n42815_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n42820_o = n41957_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n42821_o = n42820_o ? n42819_o : n42817_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n42822_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n42823_o = iregisters_r[25:13];
  assign n42824_o = iregisters_r[38:26];
  assign n42825_o = iregisters_r[51:39];
  assign n42826_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n42827_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n42828_o = iregisters_r[90:78];
  assign n42829_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n42830_o = n41961_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n42830_o)
      2'b00: n42831_o = n42822_o;
      2'b01: n42831_o = n42823_o;
      2'b10: n42831_o = n42824_o;
      2'b11: n42831_o = n42825_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n42832_o = n41961_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n42832_o)
      2'b00: n42833_o = n42826_o;
      2'b01: n42833_o = n42827_o;
      2'b10: n42833_o = n42828_o;
      2'b11: n42833_o = n42829_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n42834_o = n41961_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n42835_o = n42834_o ? n42833_o : n42831_o;
endmodule

module instr_decoder2_1_1
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n40571_o;
  wire n40573_o;
  wire n40576_o;
  wire n40578_o;
  wire n40580_o;
  wire n40582_o;
  wire [5:0] n40583_o;
  wire [3:0] n40585_o;
  wire [3:0] n40587_o;
  wire [3:0] n40588_o;
  wire [3:0] n40589_o;
  reg [3:0] n40590_o;
  wire [8:0] n40592_o;
  wire [8:0] n40594_o;
  wire [8:0] n40595_o;
  wire [8:0] n40596_o;
  reg [8:0] n40597_o;
  wire [12:0] n40600_o;
  wire n40608_o;
  wire n40610_o;
  wire n40613_o;
  wire n40615_o;
  wire n40617_o;
  wire n40619_o;
  wire [5:0] n40620_o;
  wire [3:0] n40622_o;
  wire [3:0] n40624_o;
  wire [3:0] n40625_o;
  wire [3:0] n40626_o;
  reg [3:0] n40627_o;
  wire [8:0] n40629_o;
  wire [8:0] n40631_o;
  wire [8:0] n40632_o;
  wire [8:0] n40633_o;
  reg [8:0] n40634_o;
  wire [12:0] n40637_o;
  wire [7:0] n40638_o;
  wire n40639_o;
  wire [4:0] n40640_o;
  wire [4:0] n40641_o;
  wire [11:0] n40643_o;
  wire [11:0] n40644_o;
  wire [11:0] n40645_o;
  wire [11:0] n40646_o;
  wire [3:0] n40647_o;
  wire [3:0] n40648_o;
  wire [3:0] n40649_o;
  wire [3:0] n40650_o;
  wire n40651_o;
  wire n40652_o;
  wire n40653_o;
  wire n40654_o;
  wire n40657_o;
  wire n40658_o;
  wire n40659_o;
  wire n40660_o;
  wire n40661_o;
  wire n40665_o;
  wire n40666_o;
  wire n40667_o;
  wire n40668_o;
  wire n40669_o;
  wire n40673_o;
  wire n40674_o;
  wire [51:0] n40676_o;
  wire [51:0] n40677_o;
  wire [1:0] n40678_o;
  wire n40682_o;
  wire n40683_o;
  wire n40684_o;
  wire n40685_o;
  wire [12:0] n40686_o;
  wire [1:0] n40688_o;
  wire n40692_o;
  wire n40693_o;
  wire n40694_o;
  wire n40695_o;
  wire [12:0] n40696_o;
  wire [1:0] n40698_o;
  wire n40702_o;
  wire n40703_o;
  wire n40704_o;
  wire n40705_o;
  wire [12:0] n40706_o;
  wire [1:0] n40708_o;
  wire [1:0] n40712_o;
  wire [1:0] n40717_o;
  wire [1:0] n40725_o;
  wire n40729_o;
  wire n40730_o;
  wire n40731_o;
  wire n40732_o;
  wire [12:0] n40733_o;
  wire [1:0] n40735_o;
  wire n40739_o;
  wire n40740_o;
  wire [12:0] n40741_o;
  wire n40742_o;
  wire [7:0] n40743_o;
  wire [7:0] n40744_o;
  wire n40747_o;
  wire [51:0] n40749_o;
  wire [25:0] n40750_o;
  wire n40751_o;
  wire n40752_o;
  wire [12:0] n40753_o;
  wire [12:0] n40754_o;
  wire [12:0] n40755_o;
  wire n40756_o;
  wire n40757_o;
  wire [12:0] n40758_o;
  wire [12:0] n40759_o;
  wire [12:0] n40760_o;
  wire [103:0] n40771_o;
  wire [4:0] n40796_o;
  wire [3:0] n40797_o;
  wire [3:0] n40798_o;
  wire [3:0] n40799_o;
  wire [12:0] n40800_o;
  wire n40804_o;
  wire [2:0] n40806_o;
  wire [2:0] n40810_o;
  wire n40815_o;
  wire n40816_o;
  wire n40818_o;
  wire [2:0] n40819_o;
  wire [2:0] n40821_o;
  wire n40824_o;
  wire n40826_o;
  wire n40829_o;
  wire n40831_o;
  wire [2:0] n40833_o;
  wire n40835_o;
  wire n40837_o;
  wire [2:0] n40839_o;
  wire n40841_o;
  wire [4:0] n40843_o;
  wire [1:0] n40991_o;
  wire n40993_o;
  wire n40995_o;
  wire n40996_o;
  wire [2:0] n40997_o;
  wire [12:0] n41009_o;
  wire [12:0] n41010_o;
  wire [12:0] n41011_o;
  wire [9:0] n41013_o;
  wire [12:0] n41017_o;
  wire [12:0] n41018_o;
  wire [12:0] n41020_o;
  wire [9:0] n41022_o;
  wire [12:0] n41026_o;
  wire [12:0] n41027_o;
  wire n41029_o;
  wire [1:0] n41030_o;
  wire n41032_o;
  wire n41033_o;
  wire [11:0] n41034_o;
  wire [8:0] n41035_o;
  wire [8:0] n41036_o;
  wire [2:0] n41037_o;
  wire [2:0] n41038_o;
  wire [2:0] n41039_o;
  wire n41041_o;
  wire [1:0] n41042_o;
  wire n41044_o;
  wire n41045_o;
  wire n41047_o;
  wire n41048_o;
  wire n41050_o;
  wire [4:0] n41051_o;
  wire [8:0] n41052_o;
  wire [4:0] n41053_o;
  wire [5:0] n41055_o;
  wire [2:0] n41056_o;
  wire [8:0] n41057_o;
  wire [8:0] n41058_o;
  wire [2:0] n41059_o;
  wire [12:0] n41060_o;
  wire n41061_o;
  wire [11:0] n41062_o;
  wire [8:0] n41063_o;
  wire [8:0] n41064_o;
  wire [2:0] n41065_o;
  wire n41067_o;
  wire [4:0] n41068_o;
  wire [8:0] n41069_o;
  wire [4:0] n41070_o;
  wire [5:0] n41072_o;
  wire [2:0] n41073_o;
  wire [8:0] n41074_o;
  wire [8:0] n41075_o;
  wire [2:0] n41076_o;
  wire [11:0] n41077_o;
  wire [11:0] n41078_o;
  wire [11:0] n41079_o;
  wire [11:0] n41080_o;
  wire [11:0] n41081_o;
  wire [11:0] n41084_o;
  wire [11:0] n41085_o;
  wire [1:0] n41101_o;
  wire n41103_o;
  wire n41105_o;
  wire n41106_o;
  wire [2:0] n41107_o;
  wire [12:0] n41119_o;
  wire [12:0] n41120_o;
  wire [12:0] n41121_o;
  wire [9:0] n41123_o;
  wire [12:0] n41127_o;
  wire [12:0] n41128_o;
  wire [12:0] n41130_o;
  wire [9:0] n41132_o;
  wire [12:0] n41136_o;
  wire [12:0] n41137_o;
  wire n41139_o;
  wire [1:0] n41140_o;
  wire n41142_o;
  wire n41143_o;
  wire [11:0] n41144_o;
  wire [8:0] n41145_o;
  wire [8:0] n41146_o;
  wire [2:0] n41147_o;
  wire [2:0] n41148_o;
  wire [2:0] n41149_o;
  wire n41151_o;
  wire [1:0] n41152_o;
  wire n41154_o;
  wire n41155_o;
  wire n41157_o;
  wire n41158_o;
  wire n41160_o;
  wire [4:0] n41161_o;
  wire [8:0] n41162_o;
  wire [4:0] n41163_o;
  wire [5:0] n41165_o;
  wire [2:0] n41166_o;
  wire [8:0] n41167_o;
  wire [8:0] n41168_o;
  wire [2:0] n41169_o;
  wire [12:0] n41170_o;
  wire n41171_o;
  wire [11:0] n41172_o;
  wire [8:0] n41173_o;
  wire [8:0] n41174_o;
  wire [2:0] n41175_o;
  wire n41177_o;
  wire [4:0] n41178_o;
  wire [8:0] n41179_o;
  wire [4:0] n41180_o;
  wire [5:0] n41182_o;
  wire [2:0] n41183_o;
  wire [8:0] n41184_o;
  wire [8:0] n41185_o;
  wire [2:0] n41186_o;
  wire [11:0] n41187_o;
  wire [11:0] n41188_o;
  wire [11:0] n41189_o;
  wire [11:0] n41190_o;
  wire [11:0] n41191_o;
  wire [11:0] n41194_o;
  wire [11:0] n41195_o;
  wire [1:0] n41211_o;
  wire n41213_o;
  wire n41215_o;
  wire n41216_o;
  wire [2:0] n41217_o;
  wire [12:0] n41229_o;
  wire [12:0] n41230_o;
  wire [12:0] n41231_o;
  wire [9:0] n41233_o;
  wire [12:0] n41237_o;
  wire [12:0] n41238_o;
  wire [12:0] n41240_o;
  wire [9:0] n41242_o;
  wire [12:0] n41246_o;
  wire [12:0] n41247_o;
  wire n41249_o;
  wire [1:0] n41250_o;
  wire n41252_o;
  wire n41253_o;
  wire [11:0] n41254_o;
  wire [8:0] n41255_o;
  wire [8:0] n41256_o;
  wire [2:0] n41257_o;
  wire [2:0] n41258_o;
  wire [2:0] n41259_o;
  wire n41261_o;
  wire [1:0] n41262_o;
  wire n41264_o;
  wire n41265_o;
  wire n41267_o;
  wire n41268_o;
  wire n41270_o;
  wire [4:0] n41271_o;
  wire [8:0] n41272_o;
  wire [4:0] n41273_o;
  wire [5:0] n41275_o;
  wire [2:0] n41276_o;
  wire [8:0] n41277_o;
  wire [8:0] n41278_o;
  wire [2:0] n41279_o;
  wire [12:0] n41280_o;
  wire n41281_o;
  wire [11:0] n41282_o;
  wire [8:0] n41283_o;
  wire [8:0] n41284_o;
  wire [2:0] n41285_o;
  wire n41287_o;
  wire [4:0] n41288_o;
  wire [8:0] n41289_o;
  wire [4:0] n41290_o;
  wire [5:0] n41292_o;
  wire [2:0] n41293_o;
  wire [8:0] n41294_o;
  wire [8:0] n41295_o;
  wire [2:0] n41296_o;
  wire [11:0] n41297_o;
  wire [11:0] n41298_o;
  wire [11:0] n41299_o;
  wire [11:0] n41300_o;
  wire [11:0] n41301_o;
  wire [11:0] n41304_o;
  wire [11:0] n41305_o;
  wire [1:0] n41321_o;
  wire n41323_o;
  wire n41325_o;
  wire n41326_o;
  wire [2:0] n41327_o;
  wire [12:0] n41339_o;
  wire [12:0] n41340_o;
  wire [12:0] n41341_o;
  wire [9:0] n41343_o;
  wire [12:0] n41347_o;
  wire [12:0] n41348_o;
  wire [12:0] n41350_o;
  wire [9:0] n41352_o;
  wire [12:0] n41356_o;
  wire [12:0] n41357_o;
  wire n41359_o;
  wire [1:0] n41360_o;
  wire n41362_o;
  wire n41363_o;
  wire [11:0] n41364_o;
  wire [8:0] n41365_o;
  wire [8:0] n41366_o;
  wire [2:0] n41367_o;
  wire [2:0] n41368_o;
  wire [2:0] n41369_o;
  wire n41371_o;
  wire [1:0] n41372_o;
  wire n41374_o;
  wire n41375_o;
  wire n41377_o;
  wire n41378_o;
  wire n41380_o;
  wire [4:0] n41381_o;
  wire [8:0] n41382_o;
  wire [4:0] n41383_o;
  wire [5:0] n41385_o;
  wire [2:0] n41386_o;
  wire [8:0] n41387_o;
  wire [8:0] n41388_o;
  wire [2:0] n41389_o;
  wire [12:0] n41390_o;
  wire n41391_o;
  wire [11:0] n41392_o;
  wire [8:0] n41393_o;
  wire [8:0] n41394_o;
  wire [2:0] n41395_o;
  wire n41397_o;
  wire [4:0] n41398_o;
  wire [8:0] n41399_o;
  wire [4:0] n41400_o;
  wire [5:0] n41402_o;
  wire [2:0] n41403_o;
  wire [8:0] n41404_o;
  wire [8:0] n41405_o;
  wire [2:0] n41406_o;
  wire [11:0] n41407_o;
  wire [11:0] n41408_o;
  wire [11:0] n41409_o;
  wire [11:0] n41410_o;
  wire [11:0] n41411_o;
  wire [11:0] n41414_o;
  wire [11:0] n41415_o;
  wire n41422_o;
  wire [11:0] n41424_o;
  wire [6:0] n41425_o;
  wire [7:0] n41426_o;
  wire [3:0] n41428_o;
  wire [7:0] n41429_o;
  wire [6:0] n41430_o;
  wire [7:0] n41431_o;
  wire [7:0] n41432_o;
  wire n41435_o;
  wire n41437_o;
  wire n41439_o;
  wire n41441_o;
  wire n41443_o;
  wire [4:0] n41445_o;
  wire [7:0] n41450_o;
  wire [7:0] n41452_o;
  wire [7:0] n41454_o;
  wire [7:0] n41456_o;
  reg [3:0] n41527_q;
  reg [3:0] n41528_q;
  reg [3:0] n41529_q;
  reg [3:0] n41530_q;
  reg [3:0] n41531_q;
  reg [3:0] n41532_q;
  reg n41534_q;
  reg n41535_q;
  reg [12:0] n41536_q;
  reg [12:0] n41537_q;
  reg [12:0] n41538_q;
  reg n41539_q;
  reg n41540_q;
  reg n41541_q;
  reg n41542_q;
  reg n41544_q;
  reg n41545_q;
  reg n41546_q;
  reg n41547_q;
  reg n41548_q;
  reg n41549_q;
  reg [11:0] n41550_q;
  reg n41551_q;
  reg n41552_q;
  reg n41553_q;
  reg [4:0] n41554_q;
  wire [11:0] n41555_o;
  reg [11:0] n41556_q;
  wire [11:0] n41557_o;
  reg [11:0] n41558_q;
  wire [11:0] n41559_o;
  reg [11:0] n41560_q;
  reg n41561_q;
  reg n41562_q;
  reg n41563_q;
  reg n41564_q;
  reg n41565_q;
  reg n41566_q;
  reg [4:0] n41568_q;
  reg [3:0] n41569_q;
  reg [3:0] n41570_q;
  reg [3:0] n41571_q;
  reg [12:0] n41572_q;
  reg [4:0] n41573_q;
  reg [3:0] n41574_q;
  reg [3:0] n41575_q;
  reg [3:0] n41576_q;
  reg [3:0] n41577_q;
  reg [3:0] n41578_q;
  reg [12:0] n41579_q;
  reg [12:0] n41580_q;
  reg [2:0] n41581_q;
  reg [2:0] n41582_q;
  reg [2:0] n41583_q;
  reg [2:0] n41584_q;
  reg n41586_q;
  reg n41587_q;
  reg n41588_q;
  reg n41589_q;
  reg [4:0] n41591_q;
  reg [103:0] n41592_q;
  reg [12:0] n41593_q;
  reg [12:0] n41594_q;
  reg [12:0] n41595_q;
  reg [12:0] n41596_q;
  reg [12:0] n41597_q;
  reg [12:0] n41598_q;
  reg [7:0] n41599_q;
  reg [7:0] n41600_q;
  reg [7:0] n41601_q;
  reg [7:0] n41602_q;
  reg [7:0] n41603_q;
  reg [7:0] n41604_q;
  reg [7:0] n41605_q;
  reg [7:0] n41606_q;
  reg [7:0] n41607_q;
  reg [12:0] n41608_q;
  wire [12:0] n41609_o;
  wire [12:0] n41610_o;
  wire [12:0] n41611_o;
  wire [12:0] n41612_o;
  wire [1:0] n41613_o;
  reg [12:0] n41614_o;
  wire [12:0] n41615_o;
  wire [12:0] n41616_o;
  wire [12:0] n41617_o;
  wire [12:0] n41618_o;
  wire [1:0] n41619_o;
  reg [12:0] n41620_o;
  wire [12:0] n41621_o;
  wire [12:0] n41622_o;
  wire [12:0] n41623_o;
  wire [12:0] n41624_o;
  wire [1:0] n41625_o;
  reg [12:0] n41626_o;
  wire [12:0] n41627_o;
  wire [12:0] n41628_o;
  wire [12:0] n41629_o;
  wire [12:0] n41630_o;
  wire [1:0] n41631_o;
  reg [12:0] n41632_o;
  wire [12:0] n41633_o;
  wire [12:0] n41634_o;
  wire [12:0] n41635_o;
  wire [12:0] n41636_o;
  wire [1:0] n41637_o;
  reg [12:0] n41638_o;
  wire [12:0] n41639_o;
  wire [12:0] n41640_o;
  wire [12:0] n41641_o;
  wire [12:0] n41642_o;
  wire [1:0] n41643_o;
  reg [12:0] n41644_o;
  wire [12:0] n41645_o;
  wire [12:0] n41646_o;
  wire [12:0] n41647_o;
  wire [12:0] n41648_o;
  wire [1:0] n41649_o;
  reg [12:0] n41650_o;
  wire [12:0] n41651_o;
  wire [12:0] n41652_o;
  wire [12:0] n41653_o;
  wire [12:0] n41654_o;
  wire [1:0] n41655_o;
  reg [12:0] n41656_o;
  wire [12:0] n41657_o;
  wire [12:0] n41658_o;
  wire [12:0] n41659_o;
  wire [12:0] n41660_o;
  wire [12:0] n41661_o;
  wire [12:0] n41662_o;
  wire [12:0] n41663_o;
  wire [12:0] n41664_o;
  wire [1:0] n41665_o;
  reg [12:0] n41666_o;
  wire [1:0] n41667_o;
  reg [12:0] n41668_o;
  wire n41669_o;
  wire [12:0] n41670_o;
  wire [12:0] n41671_o;
  wire [12:0] n41672_o;
  wire [12:0] n41673_o;
  wire [12:0] n41674_o;
  wire [12:0] n41675_o;
  wire [12:0] n41676_o;
  wire [12:0] n41677_o;
  wire [12:0] n41678_o;
  wire [1:0] n41679_o;
  reg [12:0] n41680_o;
  wire [1:0] n41681_o;
  reg [12:0] n41682_o;
  wire n41683_o;
  wire [12:0] n41684_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n40743_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n40600_o;
  assign i_x2_out = n40637_o;
  assign result_waddr_out = n40638_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n41527_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n41528_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n41529_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n41530_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n41531_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n41532_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n41534_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n41535_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n41536_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n41537_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n41538_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n41539_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n41540_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n41541_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n41542_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n40641_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n41544_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n41545_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n40639_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n41546_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n40661_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n41547_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n40669_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n41548_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n40674_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n41549_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n41550_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n40643_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n40644_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n40645_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n40646_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n40647_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n40648_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n40649_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n40650_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n40651_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n40652_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n40653_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n40654_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n41551_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n41552_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n41553_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n41554_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n41556_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n41558_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n41560_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n41085_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n41195_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n41305_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n41415_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n41561_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n41562_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n41563_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n41564_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n41565_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n41566_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n40796_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n40797_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n40798_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n40799_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n40800_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n41568_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n41569_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n41570_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n41571_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n41572_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n41573_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n41574_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n41575_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n41576_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n41577_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n41578_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n41579_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n41580_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n41581_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n41582_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n41583_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n41584_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n41586_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n41587_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n41588_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n41589_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n41591_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n41592_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n40676_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n40677_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n41593_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n41594_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n41595_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n41596_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n41597_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n41598_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n40686_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n40696_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n40706_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n41632_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n41638_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n41644_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n40741_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n40733_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n41656_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n41599_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n41600_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n41601_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n41602_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n41603_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n41604_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n41605_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n41606_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n41607_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n41608_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n40571_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n40573_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n40576_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n40578_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n40580_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n40582_o = imu_x1_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40583_o = {n40582_o, n40580_o, n40578_o, n40576_o, n40573_o, n40571_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40585_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40587_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40588_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40589_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n40583_o)
      6'b100000: n40590_o = n40588_o;
      6'b010000: n40590_o = n40587_o;
      6'b001000: n40590_o = 4'b0101;
      6'b000100: n40590_o = instruction_tid_rrr;
      6'b000010: n40590_o = n40585_o;
      6'b000001: n40590_o = 4'b0000;
      default: n40590_o = n40589_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40592_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40594_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40595_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40596_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n40583_o)
      6'b100000: n40597_o = n40595_o;
      6'b010000: n40597_o = n40594_o;
      6'b001000: n40597_o = 9'b000000000;
      6'b000100: n40597_o = 9'b000000000;
      6'b000010: n40597_o = n40592_o;
      6'b000001: n40597_o = 9'b000000000;
      default: n40597_o = n40596_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40600_o = {n40597_o, n40590_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n40608_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n40610_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n40613_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n40615_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n40617_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n40619_o = imu_x2_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40620_o = {n40619_o, n40617_o, n40615_o, n40613_o, n40610_o, n40608_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40622_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40624_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40625_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n40626_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n40620_o)
      6'b100000: n40627_o = n40625_o;
      6'b010000: n40627_o = n40624_o;
      6'b001000: n40627_o = 4'b0101;
      6'b000100: n40627_o = instruction_tid_rrr;
      6'b000010: n40627_o = n40622_o;
      6'b000001: n40627_o = 4'b0000;
      default: n40627_o = n40626_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40629_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40631_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40632_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40633_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n40620_o)
      6'b100000: n40634_o = n40632_o;
      6'b010000: n40634_o = n40631_o;
      6'b001000: n40634_o = 9'b000000000;
      6'b000100: n40634_o = 9'b000000000;
      6'b000010: n40634_o = n40629_o;
      6'b000001: n40634_o = 9'b000000000;
      default: n40634_o = n40633_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n40637_o = {n40634_o, n40627_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n40638_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n40639_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n40640_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n40641_o = instruction_mu_valid_in ? n40640_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n40643_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n40644_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n40645_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n40646_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n40647_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n40648_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n40649_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n40650_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n40651_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n40652_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n40653_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n40654_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n40657_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n40658_o = n40657_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n40659_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n40660_o = n40659_o & n40658_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n40661_o = n40660_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n40665_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n40666_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n40667_o = n40666_o & n40665_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n40668_o = n40667_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n40669_o = n40668_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n40673_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n40674_o = n40673_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n40676_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n40677_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n40678_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n40682_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n40683_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n40684_o = ~n40683_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n40685_o = n40682_o | n40684_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n40686_o = n40685_o ? n41614_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n40688_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n40692_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n40693_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n40694_o = ~n40693_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n40695_o = n40692_o | n40694_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n40696_o = n40695_o ? n41620_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n40698_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n40702_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n40703_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n40704_o = ~n40703_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n40705_o = n40702_o | n40704_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n40706_o = n40705_o ? n41626_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n40708_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n40712_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n40717_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n40725_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n40729_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n40730_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n40731_o = ~n40730_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n40732_o = n40729_o | n40731_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n40733_o = n40732_o ? n41650_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n40735_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n40739_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n40740_o = ~n40739_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n40741_o = n40740_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n40742_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n40743_o = n40742_o ? mu_lane_rrrrrr : n40744_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n40744_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n40747_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n40749_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n40750_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n40751_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n40752_o = ~n40751_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n40753_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n40754_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n40755_o = n40752_o ? n40753_o : n40754_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n40756_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n40757_o = ~n40756_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n40758_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n40759_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n40760_o = n40757_o ? n40758_o : n40759_o;
  assign n40771_o = {n40749_o, n40755_o, n40760_o, n40750_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n40796_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n40797_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n40798_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n40799_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n40800_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n40804_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n40806_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n40810_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n40815_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n40816_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n40818_o = n40816_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n40819_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n40821_o = n40818_o ? n40819_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n40824_o = n40818_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n40826_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n40829_o = n40826_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n40831_o = n40815_o ? n40829_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n40833_o = n40815_o ? n40821_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n40835_o = n40815_o ? n40824_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n40837_o = got_imu_rr ? n40831_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n40839_o = got_imu_rr ? n40833_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n40841_o = got_imu_rr ? n40835_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n40843_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n40991_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n40993_o = n40991_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n40995_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n40996_o = n40993_o | n40995_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n40997_o = mu_x1_parm1[2:0];
  assign n41009_o = {1'b0, mu_x1_parm1};
  assign n41010_o = {10'b0000000000, n40997_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n41011_o = n40996_o ? n41010_o : n41009_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n41013_o = mu_x1_i1_1[9:0];
  assign n41017_o = {n41013_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n41018_o = mu_x1_vector ? n41017_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n41020_o = mu_x1_i0_1 + n41011_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n41022_o = n41020_o[9:0];
  assign n41026_o = {n41022_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41027_o = mu_x1_vector ? n41026_o : n41020_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n41029_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n41030_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n41032_o = n41030_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n41033_o = n41029_o | n41032_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n41034_o = n41027_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n41035_o = n41034_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n41036_o = ~n41035_o;
  assign n41037_o = n41026_o[2:0];
  assign n41038_o = n41020_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41039_o = mu_x1_vector ? n41037_o : n41038_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n41041_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n41042_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n41044_o = n41042_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n41045_o = n41041_o | n41044_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n41047_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n41048_o = n41045_o | n41047_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n41050_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n41051_o = n41027_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n41052_o = {n41051_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n41053_o = n41027_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n41055_o = {1'b0, n41053_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n41056_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n41057_o = {n41055_o, n41056_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n41058_o = n41050_o ? n41052_o : n41057_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n41059_o = n41027_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n41060_o = n41018_o + n41027_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n41061_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n41062_o = n41060_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n41063_o = n41062_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n41064_o = ~n41063_o;
  assign n41065_o = n41060_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n41067_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n41068_o = n41060_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n41069_o = {n41068_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n41070_o = n41060_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n41072_o = {1'b0, n41070_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n41073_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n41074_o = {n41072_o, n41073_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n41075_o = n41067_o ? n41069_o : n41074_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n41076_o = n41060_o[2:0];
  assign n41077_o = {n41075_o, n41076_o};
  assign n41078_o = {n41064_o, n41065_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n41079_o = n41061_o ? n41078_o : n41077_o;
  assign n41080_o = {n41058_o, n41059_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n41081_o = n41048_o ? n41080_o : n41079_o;
  assign n41084_o = {n41036_o, n41039_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n41085_o = n41033_o ? n41084_o : n41081_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n41101_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n41103_o = n41101_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n41105_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n41106_o = n41103_o | n41105_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n41107_o = mu_x2_parm1[2:0];
  assign n41119_o = {1'b0, mu_x2_parm1};
  assign n41120_o = {10'b0000000000, n41107_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n41121_o = n41106_o ? n41120_o : n41119_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n41123_o = mu_x2_i1_1[9:0];
  assign n41127_o = {n41123_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n41128_o = mu_x2_vector ? n41127_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n41130_o = mu_x2_i0_1 + n41121_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n41132_o = n41130_o[9:0];
  assign n41136_o = {n41132_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41137_o = mu_x2_vector ? n41136_o : n41130_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n41139_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n41140_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n41142_o = n41140_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n41143_o = n41139_o | n41142_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n41144_o = n41137_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n41145_o = n41144_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n41146_o = ~n41145_o;
  assign n41147_o = n41136_o[2:0];
  assign n41148_o = n41130_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41149_o = mu_x2_vector ? n41147_o : n41148_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n41151_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n41152_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n41154_o = n41152_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n41155_o = n41151_o | n41154_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n41157_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n41158_o = n41155_o | n41157_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n41160_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n41161_o = n41137_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n41162_o = {n41161_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n41163_o = n41137_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n41165_o = {1'b0, n41163_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n41166_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n41167_o = {n41165_o, n41166_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n41168_o = n41160_o ? n41162_o : n41167_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n41169_o = n41137_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n41170_o = n41128_o + n41137_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n41171_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n41172_o = n41170_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n41173_o = n41172_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n41174_o = ~n41173_o;
  assign n41175_o = n41170_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n41177_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n41178_o = n41170_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n41179_o = {n41178_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n41180_o = n41170_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n41182_o = {1'b0, n41180_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n41183_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n41184_o = {n41182_o, n41183_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n41185_o = n41177_o ? n41179_o : n41184_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n41186_o = n41170_o[2:0];
  assign n41187_o = {n41185_o, n41186_o};
  assign n41188_o = {n41174_o, n41175_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n41189_o = n41171_o ? n41188_o : n41187_o;
  assign n41190_o = {n41168_o, n41169_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n41191_o = n41158_o ? n41190_o : n41189_o;
  assign n41194_o = {n41146_o, n41149_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n41195_o = n41143_o ? n41194_o : n41191_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n41211_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n41213_o = n41211_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n41215_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n41216_o = n41213_o | n41215_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n41217_o = mu_x3_parm1[2:0];
  assign n41229_o = {1'b0, mu_x3_parm1};
  assign n41230_o = {10'b0000000000, n41217_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n41231_o = n41216_o ? n41230_o : n41229_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n41233_o = mu_x3_i1_1[9:0];
  assign n41237_o = {n41233_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n41238_o = mu_x3_vector ? n41237_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n41240_o = mu_x3_i0_1 + n41231_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n41242_o = n41240_o[9:0];
  assign n41246_o = {n41242_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41247_o = mu_x3_vector ? n41246_o : n41240_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n41249_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n41250_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n41252_o = n41250_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n41253_o = n41249_o | n41252_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n41254_o = n41247_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n41255_o = n41254_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n41256_o = ~n41255_o;
  assign n41257_o = n41246_o[2:0];
  assign n41258_o = n41240_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41259_o = mu_x3_vector ? n41257_o : n41258_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n41261_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n41262_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n41264_o = n41262_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n41265_o = n41261_o | n41264_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n41267_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n41268_o = n41265_o | n41267_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n41270_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n41271_o = n41247_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n41272_o = {n41271_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n41273_o = n41247_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n41275_o = {1'b0, n41273_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n41276_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n41277_o = {n41275_o, n41276_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n41278_o = n41270_o ? n41272_o : n41277_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n41279_o = n41247_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n41280_o = n41238_o + n41247_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n41281_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n41282_o = n41280_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n41283_o = n41282_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n41284_o = ~n41283_o;
  assign n41285_o = n41280_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n41287_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n41288_o = n41280_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n41289_o = {n41288_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n41290_o = n41280_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n41292_o = {1'b0, n41290_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n41293_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n41294_o = {n41292_o, n41293_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n41295_o = n41287_o ? n41289_o : n41294_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n41296_o = n41280_o[2:0];
  assign n41297_o = {n41295_o, n41296_o};
  assign n41298_o = {n41284_o, n41285_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n41299_o = n41281_o ? n41298_o : n41297_o;
  assign n41300_o = {n41278_o, n41279_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n41301_o = n41268_o ? n41300_o : n41299_o;
  assign n41304_o = {n41256_o, n41259_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n41305_o = n41253_o ? n41304_o : n41301_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n41321_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n41323_o = n41321_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n41325_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n41326_o = n41323_o | n41325_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n41327_o = mu_y_parm1[2:0];
  assign n41339_o = {1'b0, mu_y_parm1};
  assign n41340_o = {10'b0000000000, n41327_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n41341_o = n41326_o ? n41340_o : n41339_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n41343_o = mu_y_i1_1[9:0];
  assign n41347_o = {n41343_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n41348_o = mu_y_vector ? n41347_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n41350_o = mu_y_i0_1 + n41341_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n41352_o = n41350_o[9:0];
  assign n41356_o = {n41352_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41357_o = mu_y_vector ? n41356_o : n41350_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n41359_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n41360_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n41362_o = n41360_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n41363_o = n41359_o | n41362_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n41364_o = n41357_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n41365_o = n41364_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n41366_o = ~n41365_o;
  assign n41367_o = n41356_o[2:0];
  assign n41368_o = n41350_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n41369_o = mu_y_vector ? n41367_o : n41368_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n41371_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n41372_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n41374_o = n41372_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n41375_o = n41371_o | n41374_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n41377_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n41378_o = n41375_o | n41377_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n41380_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n41381_o = n41357_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n41382_o = {n41381_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n41383_o = n41357_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n41385_o = {1'b0, n41383_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n41386_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n41387_o = {n41385_o, n41386_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n41388_o = n41380_o ? n41382_o : n41387_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n41389_o = n41357_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n41390_o = n41348_o + n41357_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n41391_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n41392_o = n41390_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n41393_o = n41392_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n41394_o = ~n41393_o;
  assign n41395_o = n41390_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n41397_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n41398_o = n41390_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n41399_o = {n41398_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n41400_o = n41390_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n41402_o = {1'b0, n41400_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n41403_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n41404_o = {n41402_o, n41403_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n41405_o = n41397_o ? n41399_o : n41404_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n41406_o = n41390_o[2:0];
  assign n41407_o = {n41405_o, n41406_o};
  assign n41408_o = {n41394_o, n41395_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n41409_o = n41391_o ? n41408_o : n41407_o;
  assign n41410_o = {n41388_o, n41389_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n41411_o = n41378_o ? n41410_o : n41409_o;
  assign n41414_o = {n41366_o, n41369_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n41415_o = n41363_o ? n41414_o : n41411_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n41422_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n41424_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n41425_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n41426_o = {instruction_vm_in, n41425_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n41428_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n41429_o = {n41428_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n41430_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n41431_o = {instruction_vm_in, n41430_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n41432_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41435_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41437_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41439_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41441_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41443_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41445_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41450_o = instruction_tid_valid_in ? n41432_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41452_o = instruction_tid_valid_in ? n41431_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41454_o = instruction_tid_valid_in ? n41429_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n41456_o = instruction_tid_valid_in ? n41426_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41527_q <= 4'b0000;
    else
      n41527_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41528_q <= 4'b0000;
    else
      n41528_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41529_q <= 4'b0000;
    else
      n41529_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41530_q <= 4'b0000;
    else
      n41530_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41531_q <= 4'b0000;
    else
      n41531_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41532_q <= 4'b0000;
    else
      n41532_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41534_q <= 1'b0;
    else
      n41534_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41535_q <= 1'b0;
    else
      n41535_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41536_q <= 13'b0000000000000;
    else
      n41536_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41537_q <= 13'b0000000000000;
    else
      n41537_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41538_q <= 13'b0000000000000;
    else
      n41538_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41539_q <= 1'b0;
    else
      n41539_q <= n40837_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41540_q <= 1'b0;
    else
      n41540_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41541_q <= 1'b0;
    else
      n41541_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41542_q <= 1'b0;
    else
      n41542_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41544_q <= 1'b0;
    else
      n41544_q <= n41435_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41545_q <= 1'b0;
    else
      n41545_q <= n41437_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41546_q <= 1'b0;
    else
      n41546_q <= n41439_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41547_q <= 1'b0;
    else
      n41547_q <= n41441_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41548_q <= 1'b0;
    else
      n41548_q <= n41443_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41549_q <= 1'b0;
    else
      n41549_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41550_q <= 12'b000000000000;
    else
      n41550_q <= n41424_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41551_q <= 1'b0;
    else
      n41551_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41552_q <= 1'b0;
    else
      n41552_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41553_q <= 1'b0;
    else
      n41553_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41554_q <= 5'b00000;
    else
      n41554_q <= n41445_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n41555_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41556_q <= 12'b000000000000;
    else
      n41556_q <= n41555_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n41557_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41558_q <= 12'b000000000000;
    else
      n41558_q <= n41557_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n41559_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41560_q <= 12'b000000000000;
    else
      n41560_q <= n41559_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41561_q <= 1'b0;
    else
      n41561_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41562_q <= 1'b0;
    else
      n41562_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41563_q <= 1'b0;
    else
      n41563_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41564_q <= 1'b0;
    else
      n41564_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41565_q <= 1'b0;
    else
      n41565_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41566_q <= 1'b0;
    else
      n41566_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41568_q <= 5'b00000;
    else
      n41568_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41569_q <= 4'b0000;
    else
      n41569_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41570_q <= 4'b0000;
    else
      n41570_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41571_q <= 4'b0000;
    else
      n41571_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41572_q <= 13'b0000000000000;
    else
      n41572_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41573_q <= 5'b00000;
    else
      n41573_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41574_q <= 4'b0000;
    else
      n41574_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41575_q <= 4'b0000;
    else
      n41575_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41576_q <= 4'b0000;
    else
      n41576_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41577_q <= 4'b0000;
    else
      n41577_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41578_q <= 4'b0000;
    else
      n41578_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41579_q <= 13'b0000000000000;
    else
      n41579_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41580_q <= 13'b0000000000000;
    else
      n41580_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41581_q <= 3'b000;
    else
      n41581_q <= n40839_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41582_q <= 3'b000;
    else
      n41582_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41583_q <= 3'b000;
    else
      n41583_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41584_q <= 3'b000;
    else
      n41584_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41586_q <= 1'b0;
    else
      n41586_q <= n40841_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41587_q <= 1'b0;
    else
      n41587_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41588_q <= 1'b0;
    else
      n41588_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41589_q <= 1'b0;
    else
      n41589_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41591_q <= 5'b00000;
    else
      n41591_q <= n40843_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n40747_o)
    if (n40747_o)
      n41592_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n41592_q <= n40771_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41593_q <= 13'b0000000000000;
    else
      n41593_q <= n41670_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41594_q <= 13'b0000000000000;
    else
      n41594_q <= n41684_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41595_q <= 13'b0000000000000;
    else
      n41595_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41596_q <= 13'b0000000000000;
    else
      n41596_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41597_q <= 13'b0000000000000;
    else
      n41597_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41598_q <= 13'b0000000000000;
    else
      n41598_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41599_q <= 8'b00000000;
    else
      n41599_q <= n41450_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41600_q <= 8'b00000000;
    else
      n41600_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41601_q <= 8'b00000000;
    else
      n41601_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41602_q <= 8'b00000000;
    else
      n41602_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41603_q <= 8'b00000000;
    else
      n41603_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41604_q <= 8'b00000000;
    else
      n41604_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41605_q <= 8'b00000000;
    else
      n41605_q <= n41452_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41606_q <= 8'b00000000;
    else
      n41606_q <= n41454_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n41422_o)
    if (n41422_o)
      n41607_q <= 8'b00000000;
    else
      n41607_q <= n41456_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n40804_o)
    if (n40804_o)
      n41608_q <= 13'b0000000000000;
    else
      n41608_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n41609_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n41610_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n41611_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n41612_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n41613_o = n40678_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n41613_o)
      2'b00: n41614_o = n41609_o;
      2'b01: n41614_o = n41610_o;
      2'b10: n41614_o = n41611_o;
      2'b11: n41614_o = n41612_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n41615_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n41616_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n41617_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n41618_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n41619_o = n40688_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n41619_o)
      2'b00: n41620_o = n41615_o;
      2'b01: n41620_o = n41616_o;
      2'b10: n41620_o = n41617_o;
      2'b11: n41620_o = n41618_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n41621_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n41622_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n41623_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n41624_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n41625_o = n40698_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n41625_o)
      2'b00: n41626_o = n41621_o;
      2'b01: n41626_o = n41622_o;
      2'b10: n41626_o = n41623_o;
      2'b11: n41626_o = n41624_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n41627_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n41628_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n41629_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n41630_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n41631_o = n40708_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n41631_o)
      2'b00: n41632_o = n41627_o;
      2'b01: n41632_o = n41628_o;
      2'b10: n41632_o = n41629_o;
      2'b11: n41632_o = n41630_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n41633_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n41634_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n41635_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n41636_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n41637_o = n40712_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n41637_o)
      2'b00: n41638_o = n41633_o;
      2'b01: n41638_o = n41634_o;
      2'b10: n41638_o = n41635_o;
      2'b11: n41638_o = n41636_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n41639_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n41640_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n41641_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n41642_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n41643_o = n40717_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n41643_o)
      2'b00: n41644_o = n41639_o;
      2'b01: n41644_o = n41640_o;
      2'b10: n41644_o = n41641_o;
      2'b11: n41644_o = n41642_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n41645_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n41646_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n41647_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n41648_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n41649_o = n40725_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n41649_o)
      2'b00: n41650_o = n41645_o;
      2'b01: n41650_o = n41646_o;
      2'b10: n41650_o = n41647_o;
      2'b11: n41650_o = n41648_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n41651_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n41652_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n41653_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n41654_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n41655_o = n40735_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n41655_o)
      2'b00: n41656_o = n41651_o;
      2'b01: n41656_o = n41652_o;
      2'b10: n41656_o = n41653_o;
      2'b11: n41656_o = n41654_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n41657_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n41658_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n41659_o = iregisters_r[38:26];
  assign n41660_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n41661_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n41662_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n41663_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n41664_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n41665_o = n40806_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n41665_o)
      2'b00: n41666_o = n41657_o;
      2'b01: n41666_o = n41658_o;
      2'b10: n41666_o = n41659_o;
      2'b11: n41666_o = n41660_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n41667_o = n40806_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n41667_o)
      2'b00: n41668_o = n41661_o;
      2'b01: n41668_o = n41662_o;
      2'b10: n41668_o = n41663_o;
      2'b11: n41668_o = n41664_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n41669_o = n40806_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n41670_o = n41669_o ? n41668_o : n41666_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n41671_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n41672_o = iregisters_r[25:13];
  assign n41673_o = iregisters_r[38:26];
  assign n41674_o = iregisters_r[51:39];
  assign n41675_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n41676_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n41677_o = iregisters_r[90:78];
  assign n41678_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n41679_o = n40810_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n41679_o)
      2'b00: n41680_o = n41671_o;
      2'b01: n41680_o = n41672_o;
      2'b10: n41680_o = n41673_o;
      2'b11: n41680_o = n41674_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n41681_o = n40810_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n41681_o)
      2'b00: n41682_o = n41675_o;
      2'b01: n41682_o = n41676_o;
      2'b10: n41682_o = n41677_o;
      2'b11: n41682_o = n41678_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n41683_o = n40810_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n41684_o = n41683_o ? n41682_o : n41680_o;
endmodule

module instr_decoder2_1_0
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n39420_o;
  wire n39422_o;
  wire n39425_o;
  wire n39427_o;
  wire n39429_o;
  wire n39431_o;
  wire [5:0] n39432_o;
  wire [3:0] n39434_o;
  wire [3:0] n39436_o;
  wire [3:0] n39437_o;
  wire [3:0] n39438_o;
  reg [3:0] n39439_o;
  wire [8:0] n39441_o;
  wire [8:0] n39443_o;
  wire [8:0] n39444_o;
  wire [8:0] n39445_o;
  reg [8:0] n39446_o;
  wire [12:0] n39449_o;
  wire n39457_o;
  wire n39459_o;
  wire n39462_o;
  wire n39464_o;
  wire n39466_o;
  wire n39468_o;
  wire [5:0] n39469_o;
  wire [3:0] n39471_o;
  wire [3:0] n39473_o;
  wire [3:0] n39474_o;
  wire [3:0] n39475_o;
  reg [3:0] n39476_o;
  wire [8:0] n39478_o;
  wire [8:0] n39480_o;
  wire [8:0] n39481_o;
  wire [8:0] n39482_o;
  reg [8:0] n39483_o;
  wire [12:0] n39486_o;
  wire [7:0] n39487_o;
  wire n39488_o;
  wire [4:0] n39489_o;
  wire [4:0] n39490_o;
  wire [11:0] n39492_o;
  wire [11:0] n39493_o;
  wire [11:0] n39494_o;
  wire [11:0] n39495_o;
  wire [3:0] n39496_o;
  wire [3:0] n39497_o;
  wire [3:0] n39498_o;
  wire [3:0] n39499_o;
  wire n39500_o;
  wire n39501_o;
  wire n39502_o;
  wire n39503_o;
  wire n39506_o;
  wire n39507_o;
  wire n39508_o;
  wire n39509_o;
  wire n39510_o;
  wire n39514_o;
  wire n39515_o;
  wire n39516_o;
  wire n39517_o;
  wire n39518_o;
  wire n39522_o;
  wire n39523_o;
  wire [51:0] n39525_o;
  wire [51:0] n39526_o;
  wire [1:0] n39527_o;
  wire n39531_o;
  wire n39532_o;
  wire n39533_o;
  wire n39534_o;
  wire [12:0] n39535_o;
  wire [1:0] n39537_o;
  wire n39541_o;
  wire n39542_o;
  wire n39543_o;
  wire n39544_o;
  wire [12:0] n39545_o;
  wire [1:0] n39547_o;
  wire n39551_o;
  wire n39552_o;
  wire n39553_o;
  wire n39554_o;
  wire [12:0] n39555_o;
  wire [1:0] n39557_o;
  wire [1:0] n39561_o;
  wire [1:0] n39566_o;
  wire [1:0] n39574_o;
  wire n39578_o;
  wire n39579_o;
  wire n39580_o;
  wire n39581_o;
  wire [12:0] n39582_o;
  wire [1:0] n39584_o;
  wire n39588_o;
  wire n39589_o;
  wire [12:0] n39590_o;
  wire n39591_o;
  wire [7:0] n39592_o;
  wire [7:0] n39593_o;
  wire n39596_o;
  wire [51:0] n39598_o;
  wire [25:0] n39599_o;
  wire n39600_o;
  wire n39601_o;
  wire [12:0] n39602_o;
  wire [12:0] n39603_o;
  wire [12:0] n39604_o;
  wire n39605_o;
  wire n39606_o;
  wire [12:0] n39607_o;
  wire [12:0] n39608_o;
  wire [12:0] n39609_o;
  wire [103:0] n39620_o;
  wire [4:0] n39645_o;
  wire [3:0] n39646_o;
  wire [3:0] n39647_o;
  wire [3:0] n39648_o;
  wire [12:0] n39649_o;
  wire n39653_o;
  wire [2:0] n39655_o;
  wire [2:0] n39659_o;
  wire n39664_o;
  wire n39665_o;
  wire n39667_o;
  wire [2:0] n39668_o;
  wire [2:0] n39670_o;
  wire n39673_o;
  wire n39675_o;
  wire n39678_o;
  wire n39680_o;
  wire [2:0] n39682_o;
  wire n39684_o;
  wire n39686_o;
  wire [2:0] n39688_o;
  wire n39690_o;
  wire [4:0] n39692_o;
  wire [1:0] n39840_o;
  wire n39842_o;
  wire n39844_o;
  wire n39845_o;
  wire [2:0] n39846_o;
  wire [12:0] n39858_o;
  wire [12:0] n39859_o;
  wire [12:0] n39860_o;
  wire [9:0] n39862_o;
  wire [12:0] n39866_o;
  wire [12:0] n39867_o;
  wire [12:0] n39869_o;
  wire [9:0] n39871_o;
  wire [12:0] n39875_o;
  wire [12:0] n39876_o;
  wire n39878_o;
  wire [1:0] n39879_o;
  wire n39881_o;
  wire n39882_o;
  wire [11:0] n39883_o;
  wire [8:0] n39884_o;
  wire [8:0] n39885_o;
  wire [2:0] n39886_o;
  wire [2:0] n39887_o;
  wire [2:0] n39888_o;
  wire n39890_o;
  wire [1:0] n39891_o;
  wire n39893_o;
  wire n39894_o;
  wire n39896_o;
  wire n39897_o;
  wire n39899_o;
  wire [4:0] n39900_o;
  wire [8:0] n39901_o;
  wire [4:0] n39902_o;
  wire [5:0] n39904_o;
  wire [2:0] n39905_o;
  wire [8:0] n39906_o;
  wire [8:0] n39907_o;
  wire [2:0] n39908_o;
  wire [12:0] n39909_o;
  wire n39910_o;
  wire [11:0] n39911_o;
  wire [8:0] n39912_o;
  wire [8:0] n39913_o;
  wire [2:0] n39914_o;
  wire n39916_o;
  wire [4:0] n39917_o;
  wire [8:0] n39918_o;
  wire [4:0] n39919_o;
  wire [5:0] n39921_o;
  wire [2:0] n39922_o;
  wire [8:0] n39923_o;
  wire [8:0] n39924_o;
  wire [2:0] n39925_o;
  wire [11:0] n39926_o;
  wire [11:0] n39927_o;
  wire [11:0] n39928_o;
  wire [11:0] n39929_o;
  wire [11:0] n39930_o;
  wire [11:0] n39933_o;
  wire [11:0] n39934_o;
  wire [1:0] n39950_o;
  wire n39952_o;
  wire n39954_o;
  wire n39955_o;
  wire [2:0] n39956_o;
  wire [12:0] n39968_o;
  wire [12:0] n39969_o;
  wire [12:0] n39970_o;
  wire [9:0] n39972_o;
  wire [12:0] n39976_o;
  wire [12:0] n39977_o;
  wire [12:0] n39979_o;
  wire [9:0] n39981_o;
  wire [12:0] n39985_o;
  wire [12:0] n39986_o;
  wire n39988_o;
  wire [1:0] n39989_o;
  wire n39991_o;
  wire n39992_o;
  wire [11:0] n39993_o;
  wire [8:0] n39994_o;
  wire [8:0] n39995_o;
  wire [2:0] n39996_o;
  wire [2:0] n39997_o;
  wire [2:0] n39998_o;
  wire n40000_o;
  wire [1:0] n40001_o;
  wire n40003_o;
  wire n40004_o;
  wire n40006_o;
  wire n40007_o;
  wire n40009_o;
  wire [4:0] n40010_o;
  wire [8:0] n40011_o;
  wire [4:0] n40012_o;
  wire [5:0] n40014_o;
  wire [2:0] n40015_o;
  wire [8:0] n40016_o;
  wire [8:0] n40017_o;
  wire [2:0] n40018_o;
  wire [12:0] n40019_o;
  wire n40020_o;
  wire [11:0] n40021_o;
  wire [8:0] n40022_o;
  wire [8:0] n40023_o;
  wire [2:0] n40024_o;
  wire n40026_o;
  wire [4:0] n40027_o;
  wire [8:0] n40028_o;
  wire [4:0] n40029_o;
  wire [5:0] n40031_o;
  wire [2:0] n40032_o;
  wire [8:0] n40033_o;
  wire [8:0] n40034_o;
  wire [2:0] n40035_o;
  wire [11:0] n40036_o;
  wire [11:0] n40037_o;
  wire [11:0] n40038_o;
  wire [11:0] n40039_o;
  wire [11:0] n40040_o;
  wire [11:0] n40043_o;
  wire [11:0] n40044_o;
  wire [1:0] n40060_o;
  wire n40062_o;
  wire n40064_o;
  wire n40065_o;
  wire [2:0] n40066_o;
  wire [12:0] n40078_o;
  wire [12:0] n40079_o;
  wire [12:0] n40080_o;
  wire [9:0] n40082_o;
  wire [12:0] n40086_o;
  wire [12:0] n40087_o;
  wire [12:0] n40089_o;
  wire [9:0] n40091_o;
  wire [12:0] n40095_o;
  wire [12:0] n40096_o;
  wire n40098_o;
  wire [1:0] n40099_o;
  wire n40101_o;
  wire n40102_o;
  wire [11:0] n40103_o;
  wire [8:0] n40104_o;
  wire [8:0] n40105_o;
  wire [2:0] n40106_o;
  wire [2:0] n40107_o;
  wire [2:0] n40108_o;
  wire n40110_o;
  wire [1:0] n40111_o;
  wire n40113_o;
  wire n40114_o;
  wire n40116_o;
  wire n40117_o;
  wire n40119_o;
  wire [4:0] n40120_o;
  wire [8:0] n40121_o;
  wire [4:0] n40122_o;
  wire [5:0] n40124_o;
  wire [2:0] n40125_o;
  wire [8:0] n40126_o;
  wire [8:0] n40127_o;
  wire [2:0] n40128_o;
  wire [12:0] n40129_o;
  wire n40130_o;
  wire [11:0] n40131_o;
  wire [8:0] n40132_o;
  wire [8:0] n40133_o;
  wire [2:0] n40134_o;
  wire n40136_o;
  wire [4:0] n40137_o;
  wire [8:0] n40138_o;
  wire [4:0] n40139_o;
  wire [5:0] n40141_o;
  wire [2:0] n40142_o;
  wire [8:0] n40143_o;
  wire [8:0] n40144_o;
  wire [2:0] n40145_o;
  wire [11:0] n40146_o;
  wire [11:0] n40147_o;
  wire [11:0] n40148_o;
  wire [11:0] n40149_o;
  wire [11:0] n40150_o;
  wire [11:0] n40153_o;
  wire [11:0] n40154_o;
  wire [1:0] n40170_o;
  wire n40172_o;
  wire n40174_o;
  wire n40175_o;
  wire [2:0] n40176_o;
  wire [12:0] n40188_o;
  wire [12:0] n40189_o;
  wire [12:0] n40190_o;
  wire [9:0] n40192_o;
  wire [12:0] n40196_o;
  wire [12:0] n40197_o;
  wire [12:0] n40199_o;
  wire [9:0] n40201_o;
  wire [12:0] n40205_o;
  wire [12:0] n40206_o;
  wire n40208_o;
  wire [1:0] n40209_o;
  wire n40211_o;
  wire n40212_o;
  wire [11:0] n40213_o;
  wire [8:0] n40214_o;
  wire [8:0] n40215_o;
  wire [2:0] n40216_o;
  wire [2:0] n40217_o;
  wire [2:0] n40218_o;
  wire n40220_o;
  wire [1:0] n40221_o;
  wire n40223_o;
  wire n40224_o;
  wire n40226_o;
  wire n40227_o;
  wire n40229_o;
  wire [4:0] n40230_o;
  wire [8:0] n40231_o;
  wire [4:0] n40232_o;
  wire [5:0] n40234_o;
  wire [2:0] n40235_o;
  wire [8:0] n40236_o;
  wire [8:0] n40237_o;
  wire [2:0] n40238_o;
  wire [12:0] n40239_o;
  wire n40240_o;
  wire [11:0] n40241_o;
  wire [8:0] n40242_o;
  wire [8:0] n40243_o;
  wire [2:0] n40244_o;
  wire n40246_o;
  wire [4:0] n40247_o;
  wire [8:0] n40248_o;
  wire [4:0] n40249_o;
  wire [5:0] n40251_o;
  wire [2:0] n40252_o;
  wire [8:0] n40253_o;
  wire [8:0] n40254_o;
  wire [2:0] n40255_o;
  wire [11:0] n40256_o;
  wire [11:0] n40257_o;
  wire [11:0] n40258_o;
  wire [11:0] n40259_o;
  wire [11:0] n40260_o;
  wire [11:0] n40263_o;
  wire [11:0] n40264_o;
  wire n40271_o;
  wire [11:0] n40273_o;
  wire [6:0] n40274_o;
  wire [7:0] n40275_o;
  wire [3:0] n40277_o;
  wire [7:0] n40278_o;
  wire [6:0] n40279_o;
  wire [7:0] n40280_o;
  wire [7:0] n40281_o;
  wire n40284_o;
  wire n40286_o;
  wire n40288_o;
  wire n40290_o;
  wire n40292_o;
  wire [4:0] n40294_o;
  wire [7:0] n40299_o;
  wire [7:0] n40301_o;
  wire [7:0] n40303_o;
  wire [7:0] n40305_o;
  reg [3:0] n40376_q;
  reg [3:0] n40377_q;
  reg [3:0] n40378_q;
  reg [3:0] n40379_q;
  reg [3:0] n40380_q;
  reg [3:0] n40381_q;
  reg n40383_q;
  reg n40384_q;
  reg [12:0] n40385_q;
  reg [12:0] n40386_q;
  reg [12:0] n40387_q;
  reg n40388_q;
  reg n40389_q;
  reg n40390_q;
  reg n40391_q;
  reg n40393_q;
  reg n40394_q;
  reg n40395_q;
  reg n40396_q;
  reg n40397_q;
  reg n40398_q;
  reg [11:0] n40399_q;
  reg n40400_q;
  reg n40401_q;
  reg n40402_q;
  reg [4:0] n40403_q;
  wire [11:0] n40404_o;
  reg [11:0] n40405_q;
  wire [11:0] n40406_o;
  reg [11:0] n40407_q;
  wire [11:0] n40408_o;
  reg [11:0] n40409_q;
  reg n40410_q;
  reg n40411_q;
  reg n40412_q;
  reg n40413_q;
  reg n40414_q;
  reg n40415_q;
  reg [4:0] n40417_q;
  reg [3:0] n40418_q;
  reg [3:0] n40419_q;
  reg [3:0] n40420_q;
  reg [12:0] n40421_q;
  reg [4:0] n40422_q;
  reg [3:0] n40423_q;
  reg [3:0] n40424_q;
  reg [3:0] n40425_q;
  reg [3:0] n40426_q;
  reg [3:0] n40427_q;
  reg [12:0] n40428_q;
  reg [12:0] n40429_q;
  reg [2:0] n40430_q;
  reg [2:0] n40431_q;
  reg [2:0] n40432_q;
  reg [2:0] n40433_q;
  reg n40435_q;
  reg n40436_q;
  reg n40437_q;
  reg n40438_q;
  reg [4:0] n40440_q;
  reg [103:0] n40441_q;
  reg [12:0] n40442_q;
  reg [12:0] n40443_q;
  reg [12:0] n40444_q;
  reg [12:0] n40445_q;
  reg [12:0] n40446_q;
  reg [12:0] n40447_q;
  reg [7:0] n40448_q;
  reg [7:0] n40449_q;
  reg [7:0] n40450_q;
  reg [7:0] n40451_q;
  reg [7:0] n40452_q;
  reg [7:0] n40453_q;
  reg [7:0] n40454_q;
  reg [7:0] n40455_q;
  reg [7:0] n40456_q;
  reg [12:0] n40457_q;
  wire [12:0] n40458_o;
  wire [12:0] n40459_o;
  wire [12:0] n40460_o;
  wire [12:0] n40461_o;
  wire [1:0] n40462_o;
  reg [12:0] n40463_o;
  wire [12:0] n40464_o;
  wire [12:0] n40465_o;
  wire [12:0] n40466_o;
  wire [12:0] n40467_o;
  wire [1:0] n40468_o;
  reg [12:0] n40469_o;
  wire [12:0] n40470_o;
  wire [12:0] n40471_o;
  wire [12:0] n40472_o;
  wire [12:0] n40473_o;
  wire [1:0] n40474_o;
  reg [12:0] n40475_o;
  wire [12:0] n40476_o;
  wire [12:0] n40477_o;
  wire [12:0] n40478_o;
  wire [12:0] n40479_o;
  wire [1:0] n40480_o;
  reg [12:0] n40481_o;
  wire [12:0] n40482_o;
  wire [12:0] n40483_o;
  wire [12:0] n40484_o;
  wire [12:0] n40485_o;
  wire [1:0] n40486_o;
  reg [12:0] n40487_o;
  wire [12:0] n40488_o;
  wire [12:0] n40489_o;
  wire [12:0] n40490_o;
  wire [12:0] n40491_o;
  wire [1:0] n40492_o;
  reg [12:0] n40493_o;
  wire [12:0] n40494_o;
  wire [12:0] n40495_o;
  wire [12:0] n40496_o;
  wire [12:0] n40497_o;
  wire [1:0] n40498_o;
  reg [12:0] n40499_o;
  wire [12:0] n40500_o;
  wire [12:0] n40501_o;
  wire [12:0] n40502_o;
  wire [12:0] n40503_o;
  wire [1:0] n40504_o;
  reg [12:0] n40505_o;
  wire [12:0] n40506_o;
  wire [12:0] n40507_o;
  wire [12:0] n40508_o;
  wire [12:0] n40509_o;
  wire [12:0] n40510_o;
  wire [12:0] n40511_o;
  wire [12:0] n40512_o;
  wire [12:0] n40513_o;
  wire [1:0] n40514_o;
  reg [12:0] n40515_o;
  wire [1:0] n40516_o;
  reg [12:0] n40517_o;
  wire n40518_o;
  wire [12:0] n40519_o;
  wire [12:0] n40520_o;
  wire [12:0] n40521_o;
  wire [12:0] n40522_o;
  wire [12:0] n40523_o;
  wire [12:0] n40524_o;
  wire [12:0] n40525_o;
  wire [12:0] n40526_o;
  wire [12:0] n40527_o;
  wire [1:0] n40528_o;
  reg [12:0] n40529_o;
  wire [1:0] n40530_o;
  reg [12:0] n40531_o;
  wire n40532_o;
  wire [12:0] n40533_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n39592_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n39449_o;
  assign i_x2_out = n39486_o;
  assign result_waddr_out = n39487_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n40376_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n40377_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n40378_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n40379_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n40380_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n40381_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n40383_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n40384_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n40385_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n40386_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n40387_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n40388_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n40389_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n40390_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n40391_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n39490_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n40393_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n40394_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n39488_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n40395_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n39510_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n40396_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n39518_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n40397_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n39523_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n40398_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n40399_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n39492_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n39493_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n39494_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n39495_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n39496_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n39497_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n39498_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n39499_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n39500_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n39501_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n39502_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n39503_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n40400_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n40401_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n40402_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n40403_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n40405_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n40407_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n40409_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n39934_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n40044_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n40154_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n40264_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n40410_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n40411_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n40412_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n40413_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n40414_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n40415_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n39645_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n39646_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n39647_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n39648_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n39649_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n40417_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n40418_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n40419_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n40420_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n40421_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n40422_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n40423_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n40424_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n40425_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n40426_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n40427_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n40428_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n40429_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n40430_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n40431_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n40432_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n40433_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n40435_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n40436_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n40437_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n40438_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n40440_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n40441_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n39525_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n39526_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n40442_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n40443_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n40444_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n40445_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n40446_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n40447_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n39535_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n39545_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n39555_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n40481_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n40487_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n40493_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n39590_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n39582_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n40505_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n40448_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n40449_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n40450_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n40451_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n40452_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n40453_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n40454_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n40455_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n40456_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n40457_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n39420_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n39422_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n39425_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n39427_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n39429_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n39431_o = imu_x1_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39432_o = {n39431_o, n39429_o, n39427_o, n39425_o, n39422_o, n39420_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39434_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39436_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39437_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39438_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n39432_o)
      6'b100000: n39439_o = n39437_o;
      6'b010000: n39439_o = n39436_o;
      6'b001000: n39439_o = 4'b0100;
      6'b000100: n39439_o = instruction_tid_rrr;
      6'b000010: n39439_o = n39434_o;
      6'b000001: n39439_o = 4'b0000;
      default: n39439_o = n39438_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39441_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39443_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39444_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39445_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n39432_o)
      6'b100000: n39446_o = n39444_o;
      6'b010000: n39446_o = n39443_o;
      6'b001000: n39446_o = 9'b000000000;
      6'b000100: n39446_o = 9'b000000000;
      6'b000010: n39446_o = n39441_o;
      6'b000001: n39446_o = 9'b000000000;
      default: n39446_o = n39445_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39449_o = {n39446_o, n39439_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n39457_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n39459_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n39462_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n39464_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n39466_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n39468_o = imu_x2_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39469_o = {n39468_o, n39466_o, n39464_o, n39462_o, n39459_o, n39457_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39471_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39473_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39474_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n39475_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n39469_o)
      6'b100000: n39476_o = n39474_o;
      6'b010000: n39476_o = n39473_o;
      6'b001000: n39476_o = 4'b0100;
      6'b000100: n39476_o = instruction_tid_rrr;
      6'b000010: n39476_o = n39471_o;
      6'b000001: n39476_o = 4'b0000;
      default: n39476_o = n39475_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39478_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39480_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39481_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39482_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n39469_o)
      6'b100000: n39483_o = n39481_o;
      6'b010000: n39483_o = n39480_o;
      6'b001000: n39483_o = 9'b000000000;
      6'b000100: n39483_o = 9'b000000000;
      6'b000010: n39483_o = n39478_o;
      6'b000001: n39483_o = 9'b000000000;
      default: n39483_o = n39482_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n39486_o = {n39483_o, n39476_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n39487_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n39488_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n39489_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n39490_o = instruction_mu_valid_in ? n39489_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n39492_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n39493_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n39494_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n39495_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n39496_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n39497_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n39498_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n39499_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n39500_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n39501_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n39502_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n39503_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n39506_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n39507_o = n39506_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n39508_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n39509_o = n39508_o & n39507_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n39510_o = n39509_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n39514_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n39515_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n39516_o = n39515_o & n39514_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n39517_o = n39516_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n39518_o = n39517_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n39522_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n39523_o = n39522_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n39525_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n39526_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n39527_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n39531_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n39532_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n39533_o = ~n39532_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n39534_o = n39531_o | n39533_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n39535_o = n39534_o ? n40463_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n39537_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n39541_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n39542_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n39543_o = ~n39542_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n39544_o = n39541_o | n39543_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n39545_o = n39544_o ? n40469_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n39547_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n39551_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n39552_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n39553_o = ~n39552_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n39554_o = n39551_o | n39553_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n39555_o = n39554_o ? n40475_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n39557_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n39561_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n39566_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n39574_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n39578_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n39579_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n39580_o = ~n39579_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n39581_o = n39578_o | n39580_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n39582_o = n39581_o ? n40499_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n39584_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n39588_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n39589_o = ~n39588_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n39590_o = n39589_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n39591_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n39592_o = n39591_o ? mu_lane_rrrrrr : n39593_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n39593_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n39596_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n39598_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n39599_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n39600_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n39601_o = ~n39600_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n39602_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n39603_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n39604_o = n39601_o ? n39602_o : n39603_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n39605_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n39606_o = ~n39605_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n39607_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n39608_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n39609_o = n39606_o ? n39607_o : n39608_o;
  assign n39620_o = {n39598_o, n39604_o, n39609_o, n39599_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n39645_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n39646_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n39647_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n39648_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n39649_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n39653_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n39655_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n39659_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n39664_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n39665_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n39667_o = n39665_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n39668_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n39670_o = n39667_o ? n39668_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n39673_o = n39667_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n39675_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n39678_o = n39675_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n39680_o = n39664_o ? n39678_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n39682_o = n39664_o ? n39670_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n39684_o = n39664_o ? n39673_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n39686_o = got_imu_rr ? n39680_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n39688_o = got_imu_rr ? n39682_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n39690_o = got_imu_rr ? n39684_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n39692_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n39840_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n39842_o = n39840_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n39844_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n39845_o = n39842_o | n39844_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n39846_o = mu_x1_parm1[2:0];
  assign n39858_o = {1'b0, mu_x1_parm1};
  assign n39859_o = {10'b0000000000, n39846_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n39860_o = n39845_o ? n39859_o : n39858_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n39862_o = mu_x1_i1_1[9:0];
  assign n39866_o = {n39862_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n39867_o = mu_x1_vector ? n39866_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n39869_o = mu_x1_i0_1 + n39860_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n39871_o = n39869_o[9:0];
  assign n39875_o = {n39871_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n39876_o = mu_x1_vector ? n39875_o : n39869_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n39878_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n39879_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n39881_o = n39879_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n39882_o = n39878_o | n39881_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n39883_o = n39876_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n39884_o = n39883_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n39885_o = ~n39884_o;
  assign n39886_o = n39875_o[2:0];
  assign n39887_o = n39869_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n39888_o = mu_x1_vector ? n39886_o : n39887_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n39890_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n39891_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n39893_o = n39891_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n39894_o = n39890_o | n39893_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n39896_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n39897_o = n39894_o | n39896_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n39899_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n39900_o = n39876_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n39901_o = {n39900_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n39902_o = n39876_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n39904_o = {1'b0, n39902_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n39905_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n39906_o = {n39904_o, n39905_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n39907_o = n39899_o ? n39901_o : n39906_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n39908_o = n39876_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n39909_o = n39867_o + n39876_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n39910_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n39911_o = n39909_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n39912_o = n39911_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n39913_o = ~n39912_o;
  assign n39914_o = n39909_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n39916_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n39917_o = n39909_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n39918_o = {n39917_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n39919_o = n39909_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n39921_o = {1'b0, n39919_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n39922_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n39923_o = {n39921_o, n39922_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n39924_o = n39916_o ? n39918_o : n39923_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n39925_o = n39909_o[2:0];
  assign n39926_o = {n39924_o, n39925_o};
  assign n39927_o = {n39913_o, n39914_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n39928_o = n39910_o ? n39927_o : n39926_o;
  assign n39929_o = {n39907_o, n39908_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n39930_o = n39897_o ? n39929_o : n39928_o;
  assign n39933_o = {n39885_o, n39888_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n39934_o = n39882_o ? n39933_o : n39930_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n39950_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n39952_o = n39950_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n39954_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n39955_o = n39952_o | n39954_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n39956_o = mu_x2_parm1[2:0];
  assign n39968_o = {1'b0, mu_x2_parm1};
  assign n39969_o = {10'b0000000000, n39956_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n39970_o = n39955_o ? n39969_o : n39968_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n39972_o = mu_x2_i1_1[9:0];
  assign n39976_o = {n39972_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n39977_o = mu_x2_vector ? n39976_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n39979_o = mu_x2_i0_1 + n39970_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n39981_o = n39979_o[9:0];
  assign n39985_o = {n39981_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n39986_o = mu_x2_vector ? n39985_o : n39979_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n39988_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n39989_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n39991_o = n39989_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n39992_o = n39988_o | n39991_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n39993_o = n39986_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n39994_o = n39993_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n39995_o = ~n39994_o;
  assign n39996_o = n39985_o[2:0];
  assign n39997_o = n39979_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n39998_o = mu_x2_vector ? n39996_o : n39997_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n40000_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n40001_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n40003_o = n40001_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n40004_o = n40000_o | n40003_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n40006_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n40007_o = n40004_o | n40006_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n40009_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n40010_o = n39986_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n40011_o = {n40010_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n40012_o = n39986_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n40014_o = {1'b0, n40012_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n40015_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n40016_o = {n40014_o, n40015_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n40017_o = n40009_o ? n40011_o : n40016_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n40018_o = n39986_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n40019_o = n39977_o + n39986_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n40020_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n40021_o = n40019_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n40022_o = n40021_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n40023_o = ~n40022_o;
  assign n40024_o = n40019_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n40026_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n40027_o = n40019_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n40028_o = {n40027_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n40029_o = n40019_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n40031_o = {1'b0, n40029_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n40032_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n40033_o = {n40031_o, n40032_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n40034_o = n40026_o ? n40028_o : n40033_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n40035_o = n40019_o[2:0];
  assign n40036_o = {n40034_o, n40035_o};
  assign n40037_o = {n40023_o, n40024_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n40038_o = n40020_o ? n40037_o : n40036_o;
  assign n40039_o = {n40017_o, n40018_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n40040_o = n40007_o ? n40039_o : n40038_o;
  assign n40043_o = {n39995_o, n39998_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n40044_o = n39992_o ? n40043_o : n40040_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n40060_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n40062_o = n40060_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n40064_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n40065_o = n40062_o | n40064_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n40066_o = mu_x3_parm1[2:0];
  assign n40078_o = {1'b0, mu_x3_parm1};
  assign n40079_o = {10'b0000000000, n40066_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n40080_o = n40065_o ? n40079_o : n40078_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n40082_o = mu_x3_i1_1[9:0];
  assign n40086_o = {n40082_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n40087_o = mu_x3_vector ? n40086_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n40089_o = mu_x3_i0_1 + n40080_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n40091_o = n40089_o[9:0];
  assign n40095_o = {n40091_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n40096_o = mu_x3_vector ? n40095_o : n40089_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n40098_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n40099_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n40101_o = n40099_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n40102_o = n40098_o | n40101_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n40103_o = n40096_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n40104_o = n40103_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n40105_o = ~n40104_o;
  assign n40106_o = n40095_o[2:0];
  assign n40107_o = n40089_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n40108_o = mu_x3_vector ? n40106_o : n40107_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n40110_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n40111_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n40113_o = n40111_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n40114_o = n40110_o | n40113_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n40116_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n40117_o = n40114_o | n40116_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n40119_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n40120_o = n40096_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n40121_o = {n40120_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n40122_o = n40096_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n40124_o = {1'b0, n40122_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n40125_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n40126_o = {n40124_o, n40125_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n40127_o = n40119_o ? n40121_o : n40126_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n40128_o = n40096_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n40129_o = n40087_o + n40096_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n40130_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n40131_o = n40129_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n40132_o = n40131_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n40133_o = ~n40132_o;
  assign n40134_o = n40129_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n40136_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n40137_o = n40129_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n40138_o = {n40137_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n40139_o = n40129_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n40141_o = {1'b0, n40139_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n40142_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n40143_o = {n40141_o, n40142_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n40144_o = n40136_o ? n40138_o : n40143_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n40145_o = n40129_o[2:0];
  assign n40146_o = {n40144_o, n40145_o};
  assign n40147_o = {n40133_o, n40134_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n40148_o = n40130_o ? n40147_o : n40146_o;
  assign n40149_o = {n40127_o, n40128_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n40150_o = n40117_o ? n40149_o : n40148_o;
  assign n40153_o = {n40105_o, n40108_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n40154_o = n40102_o ? n40153_o : n40150_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n40170_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n40172_o = n40170_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n40174_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n40175_o = n40172_o | n40174_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n40176_o = mu_y_parm1[2:0];
  assign n40188_o = {1'b0, mu_y_parm1};
  assign n40189_o = {10'b0000000000, n40176_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n40190_o = n40175_o ? n40189_o : n40188_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n40192_o = mu_y_i1_1[9:0];
  assign n40196_o = {n40192_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n40197_o = mu_y_vector ? n40196_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n40199_o = mu_y_i0_1 + n40190_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n40201_o = n40199_o[9:0];
  assign n40205_o = {n40201_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n40206_o = mu_y_vector ? n40205_o : n40199_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n40208_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n40209_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n40211_o = n40209_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n40212_o = n40208_o | n40211_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n40213_o = n40206_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n40214_o = n40213_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n40215_o = ~n40214_o;
  assign n40216_o = n40205_o[2:0];
  assign n40217_o = n40199_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n40218_o = mu_y_vector ? n40216_o : n40217_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n40220_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n40221_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n40223_o = n40221_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n40224_o = n40220_o | n40223_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n40226_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n40227_o = n40224_o | n40226_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n40229_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n40230_o = n40206_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n40231_o = {n40230_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n40232_o = n40206_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n40234_o = {1'b0, n40232_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n40235_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n40236_o = {n40234_o, n40235_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n40237_o = n40229_o ? n40231_o : n40236_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n40238_o = n40206_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n40239_o = n40197_o + n40206_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n40240_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n40241_o = n40239_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n40242_o = n40241_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n40243_o = ~n40242_o;
  assign n40244_o = n40239_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n40246_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n40247_o = n40239_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n40248_o = {n40247_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n40249_o = n40239_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n40251_o = {1'b0, n40249_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n40252_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n40253_o = {n40251_o, n40252_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n40254_o = n40246_o ? n40248_o : n40253_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n40255_o = n40239_o[2:0];
  assign n40256_o = {n40254_o, n40255_o};
  assign n40257_o = {n40243_o, n40244_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n40258_o = n40240_o ? n40257_o : n40256_o;
  assign n40259_o = {n40237_o, n40238_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n40260_o = n40227_o ? n40259_o : n40258_o;
  assign n40263_o = {n40215_o, n40218_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n40264_o = n40212_o ? n40263_o : n40260_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n40271_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n40273_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n40274_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n40275_o = {instruction_vm_in, n40274_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n40277_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n40278_o = {n40277_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n40279_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n40280_o = {instruction_vm_in, n40279_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n40281_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40284_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40286_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40288_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40290_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40292_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40294_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40299_o = instruction_tid_valid_in ? n40281_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40301_o = instruction_tid_valid_in ? n40280_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40303_o = instruction_tid_valid_in ? n40278_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n40305_o = instruction_tid_valid_in ? n40275_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40376_q <= 4'b0000;
    else
      n40376_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40377_q <= 4'b0000;
    else
      n40377_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40378_q <= 4'b0000;
    else
      n40378_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40379_q <= 4'b0000;
    else
      n40379_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40380_q <= 4'b0000;
    else
      n40380_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40381_q <= 4'b0000;
    else
      n40381_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40383_q <= 1'b0;
    else
      n40383_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40384_q <= 1'b0;
    else
      n40384_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40385_q <= 13'b0000000000000;
    else
      n40385_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40386_q <= 13'b0000000000000;
    else
      n40386_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40387_q <= 13'b0000000000000;
    else
      n40387_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40388_q <= 1'b0;
    else
      n40388_q <= n39686_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40389_q <= 1'b0;
    else
      n40389_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40390_q <= 1'b0;
    else
      n40390_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40391_q <= 1'b0;
    else
      n40391_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40393_q <= 1'b0;
    else
      n40393_q <= n40284_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40394_q <= 1'b0;
    else
      n40394_q <= n40286_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40395_q <= 1'b0;
    else
      n40395_q <= n40288_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40396_q <= 1'b0;
    else
      n40396_q <= n40290_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40397_q <= 1'b0;
    else
      n40397_q <= n40292_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40398_q <= 1'b0;
    else
      n40398_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40399_q <= 12'b000000000000;
    else
      n40399_q <= n40273_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40400_q <= 1'b0;
    else
      n40400_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40401_q <= 1'b0;
    else
      n40401_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40402_q <= 1'b0;
    else
      n40402_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40403_q <= 5'b00000;
    else
      n40403_q <= n40294_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n40404_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40405_q <= 12'b000000000000;
    else
      n40405_q <= n40404_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n40406_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40407_q <= 12'b000000000000;
    else
      n40407_q <= n40406_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n40408_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40409_q <= 12'b000000000000;
    else
      n40409_q <= n40408_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40410_q <= 1'b0;
    else
      n40410_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40411_q <= 1'b0;
    else
      n40411_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40412_q <= 1'b0;
    else
      n40412_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40413_q <= 1'b0;
    else
      n40413_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40414_q <= 1'b0;
    else
      n40414_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40415_q <= 1'b0;
    else
      n40415_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40417_q <= 5'b00000;
    else
      n40417_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40418_q <= 4'b0000;
    else
      n40418_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40419_q <= 4'b0000;
    else
      n40419_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40420_q <= 4'b0000;
    else
      n40420_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40421_q <= 13'b0000000000000;
    else
      n40421_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40422_q <= 5'b00000;
    else
      n40422_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40423_q <= 4'b0000;
    else
      n40423_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40424_q <= 4'b0000;
    else
      n40424_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40425_q <= 4'b0000;
    else
      n40425_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40426_q <= 4'b0000;
    else
      n40426_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40427_q <= 4'b0000;
    else
      n40427_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40428_q <= 13'b0000000000000;
    else
      n40428_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40429_q <= 13'b0000000000000;
    else
      n40429_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40430_q <= 3'b000;
    else
      n40430_q <= n39688_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40431_q <= 3'b000;
    else
      n40431_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40432_q <= 3'b000;
    else
      n40432_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40433_q <= 3'b000;
    else
      n40433_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40435_q <= 1'b0;
    else
      n40435_q <= n39690_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40436_q <= 1'b0;
    else
      n40436_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40437_q <= 1'b0;
    else
      n40437_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40438_q <= 1'b0;
    else
      n40438_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40440_q <= 5'b00000;
    else
      n40440_q <= n39692_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n39596_o)
    if (n39596_o)
      n40441_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n40441_q <= n39620_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40442_q <= 13'b0000000000000;
    else
      n40442_q <= n40519_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40443_q <= 13'b0000000000000;
    else
      n40443_q <= n40533_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40444_q <= 13'b0000000000000;
    else
      n40444_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40445_q <= 13'b0000000000000;
    else
      n40445_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40446_q <= 13'b0000000000000;
    else
      n40446_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40447_q <= 13'b0000000000000;
    else
      n40447_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40448_q <= 8'b00000000;
    else
      n40448_q <= n40299_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40449_q <= 8'b00000000;
    else
      n40449_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40450_q <= 8'b00000000;
    else
      n40450_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40451_q <= 8'b00000000;
    else
      n40451_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40452_q <= 8'b00000000;
    else
      n40452_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40453_q <= 8'b00000000;
    else
      n40453_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40454_q <= 8'b00000000;
    else
      n40454_q <= n40301_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40455_q <= 8'b00000000;
    else
      n40455_q <= n40303_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n40271_o)
    if (n40271_o)
      n40456_q <= 8'b00000000;
    else
      n40456_q <= n40305_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n39653_o)
    if (n39653_o)
      n40457_q <= 13'b0000000000000;
    else
      n40457_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n40458_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n40459_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n40460_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n40461_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n40462_o = n39527_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n40462_o)
      2'b00: n40463_o = n40458_o;
      2'b01: n40463_o = n40459_o;
      2'b10: n40463_o = n40460_o;
      2'b11: n40463_o = n40461_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n40464_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n40465_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n40466_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n40467_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n40468_o = n39537_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n40468_o)
      2'b00: n40469_o = n40464_o;
      2'b01: n40469_o = n40465_o;
      2'b10: n40469_o = n40466_o;
      2'b11: n40469_o = n40467_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n40470_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n40471_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n40472_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n40473_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n40474_o = n39547_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n40474_o)
      2'b00: n40475_o = n40470_o;
      2'b01: n40475_o = n40471_o;
      2'b10: n40475_o = n40472_o;
      2'b11: n40475_o = n40473_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n40476_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n40477_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n40478_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n40479_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n40480_o = n39557_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n40480_o)
      2'b00: n40481_o = n40476_o;
      2'b01: n40481_o = n40477_o;
      2'b10: n40481_o = n40478_o;
      2'b11: n40481_o = n40479_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n40482_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n40483_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n40484_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n40485_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n40486_o = n39561_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n40486_o)
      2'b00: n40487_o = n40482_o;
      2'b01: n40487_o = n40483_o;
      2'b10: n40487_o = n40484_o;
      2'b11: n40487_o = n40485_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n40488_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n40489_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n40490_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n40491_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n40492_o = n39566_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n40492_o)
      2'b00: n40493_o = n40488_o;
      2'b01: n40493_o = n40489_o;
      2'b10: n40493_o = n40490_o;
      2'b11: n40493_o = n40491_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n40494_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n40495_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n40496_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n40497_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n40498_o = n39574_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n40498_o)
      2'b00: n40499_o = n40494_o;
      2'b01: n40499_o = n40495_o;
      2'b10: n40499_o = n40496_o;
      2'b11: n40499_o = n40497_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n40500_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n40501_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n40502_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n40503_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n40504_o = n39584_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n40504_o)
      2'b00: n40505_o = n40500_o;
      2'b01: n40505_o = n40501_o;
      2'b10: n40505_o = n40502_o;
      2'b11: n40505_o = n40503_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n40506_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n40507_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n40508_o = iregisters_r[38:26];
  assign n40509_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n40510_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n40511_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n40512_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n40513_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n40514_o = n39655_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n40514_o)
      2'b00: n40515_o = n40506_o;
      2'b01: n40515_o = n40507_o;
      2'b10: n40515_o = n40508_o;
      2'b11: n40515_o = n40509_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n40516_o = n39655_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n40516_o)
      2'b00: n40517_o = n40510_o;
      2'b01: n40517_o = n40511_o;
      2'b10: n40517_o = n40512_o;
      2'b11: n40517_o = n40513_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n40518_o = n39655_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n40519_o = n40518_o ? n40517_o : n40515_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n40520_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n40521_o = iregisters_r[25:13];
  assign n40522_o = iregisters_r[38:26];
  assign n40523_o = iregisters_r[51:39];
  assign n40524_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n40525_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n40526_o = iregisters_r[90:78];
  assign n40527_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n40528_o = n39659_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n40528_o)
      2'b00: n40529_o = n40520_o;
      2'b01: n40529_o = n40521_o;
      2'b10: n40529_o = n40522_o;
      2'b11: n40529_o = n40523_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n40530_o = n39659_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n40530_o)
      2'b00: n40531_o = n40524_o;
      2'b01: n40531_o = n40525_o;
      2'b10: n40531_o = n40526_o;
      2'b11: n40531_o = n40527_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n40532_o = n39659_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n40533_o = n40532_o ? n40531_o : n40529_o;
endmodule

module instr_decoder2_0_3
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n38269_o;
  wire n38271_o;
  wire n38274_o;
  wire n38276_o;
  wire n38278_o;
  wire n38280_o;
  wire [5:0] n38281_o;
  wire [3:0] n38283_o;
  wire [3:0] n38285_o;
  wire [3:0] n38286_o;
  wire [3:0] n38287_o;
  reg [3:0] n38288_o;
  wire [8:0] n38290_o;
  wire [8:0] n38292_o;
  wire [8:0] n38293_o;
  wire [8:0] n38294_o;
  reg [8:0] n38295_o;
  wire [12:0] n38298_o;
  wire n38306_o;
  wire n38308_o;
  wire n38311_o;
  wire n38313_o;
  wire n38315_o;
  wire n38317_o;
  wire [5:0] n38318_o;
  wire [3:0] n38320_o;
  wire [3:0] n38322_o;
  wire [3:0] n38323_o;
  wire [3:0] n38324_o;
  reg [3:0] n38325_o;
  wire [8:0] n38327_o;
  wire [8:0] n38329_o;
  wire [8:0] n38330_o;
  wire [8:0] n38331_o;
  reg [8:0] n38332_o;
  wire [12:0] n38335_o;
  wire [7:0] n38336_o;
  wire n38337_o;
  wire [4:0] n38338_o;
  wire [4:0] n38339_o;
  wire [11:0] n38341_o;
  wire [11:0] n38342_o;
  wire [11:0] n38343_o;
  wire [11:0] n38344_o;
  wire [3:0] n38345_o;
  wire [3:0] n38346_o;
  wire [3:0] n38347_o;
  wire [3:0] n38348_o;
  wire n38349_o;
  wire n38350_o;
  wire n38351_o;
  wire n38352_o;
  wire n38355_o;
  wire n38356_o;
  wire n38357_o;
  wire n38358_o;
  wire n38359_o;
  wire n38363_o;
  wire n38364_o;
  wire n38365_o;
  wire n38366_o;
  wire n38367_o;
  wire n38371_o;
  wire n38372_o;
  wire [51:0] n38374_o;
  wire [51:0] n38375_o;
  wire [1:0] n38376_o;
  wire n38380_o;
  wire n38381_o;
  wire n38382_o;
  wire n38383_o;
  wire [12:0] n38384_o;
  wire [1:0] n38386_o;
  wire n38390_o;
  wire n38391_o;
  wire n38392_o;
  wire n38393_o;
  wire [12:0] n38394_o;
  wire [1:0] n38396_o;
  wire n38400_o;
  wire n38401_o;
  wire n38402_o;
  wire n38403_o;
  wire [12:0] n38404_o;
  wire [1:0] n38406_o;
  wire [1:0] n38410_o;
  wire [1:0] n38415_o;
  wire [1:0] n38423_o;
  wire n38427_o;
  wire n38428_o;
  wire n38429_o;
  wire n38430_o;
  wire [12:0] n38431_o;
  wire [1:0] n38433_o;
  wire n38437_o;
  wire n38438_o;
  wire [12:0] n38439_o;
  wire n38440_o;
  wire [7:0] n38441_o;
  wire [7:0] n38442_o;
  wire n38445_o;
  wire [51:0] n38447_o;
  wire [25:0] n38448_o;
  wire n38449_o;
  wire n38450_o;
  wire [12:0] n38451_o;
  wire [12:0] n38452_o;
  wire [12:0] n38453_o;
  wire n38454_o;
  wire n38455_o;
  wire [12:0] n38456_o;
  wire [12:0] n38457_o;
  wire [12:0] n38458_o;
  wire [103:0] n38469_o;
  wire [4:0] n38494_o;
  wire [3:0] n38495_o;
  wire [3:0] n38496_o;
  wire [3:0] n38497_o;
  wire [12:0] n38498_o;
  wire n38502_o;
  wire [2:0] n38504_o;
  wire [2:0] n38508_o;
  wire n38513_o;
  wire n38514_o;
  wire n38516_o;
  wire [2:0] n38517_o;
  wire [2:0] n38519_o;
  wire n38522_o;
  wire n38524_o;
  wire n38527_o;
  wire n38529_o;
  wire [2:0] n38531_o;
  wire n38533_o;
  wire n38535_o;
  wire [2:0] n38537_o;
  wire n38539_o;
  wire [4:0] n38541_o;
  wire [1:0] n38689_o;
  wire n38691_o;
  wire n38693_o;
  wire n38694_o;
  wire [2:0] n38695_o;
  wire [12:0] n38707_o;
  wire [12:0] n38708_o;
  wire [12:0] n38709_o;
  wire [9:0] n38711_o;
  wire [12:0] n38715_o;
  wire [12:0] n38716_o;
  wire [12:0] n38718_o;
  wire [9:0] n38720_o;
  wire [12:0] n38724_o;
  wire [12:0] n38725_o;
  wire n38727_o;
  wire [1:0] n38728_o;
  wire n38730_o;
  wire n38731_o;
  wire [11:0] n38732_o;
  wire [8:0] n38733_o;
  wire [8:0] n38734_o;
  wire [2:0] n38735_o;
  wire [2:0] n38736_o;
  wire [2:0] n38737_o;
  wire n38739_o;
  wire [1:0] n38740_o;
  wire n38742_o;
  wire n38743_o;
  wire n38745_o;
  wire n38746_o;
  wire n38748_o;
  wire [4:0] n38749_o;
  wire [8:0] n38750_o;
  wire [4:0] n38751_o;
  wire [5:0] n38753_o;
  wire [2:0] n38754_o;
  wire [8:0] n38755_o;
  wire [8:0] n38756_o;
  wire [2:0] n38757_o;
  wire [12:0] n38758_o;
  wire n38759_o;
  wire [11:0] n38760_o;
  wire [8:0] n38761_o;
  wire [8:0] n38762_o;
  wire [2:0] n38763_o;
  wire n38765_o;
  wire [4:0] n38766_o;
  wire [8:0] n38767_o;
  wire [4:0] n38768_o;
  wire [5:0] n38770_o;
  wire [2:0] n38771_o;
  wire [8:0] n38772_o;
  wire [8:0] n38773_o;
  wire [2:0] n38774_o;
  wire [11:0] n38775_o;
  wire [11:0] n38776_o;
  wire [11:0] n38777_o;
  wire [11:0] n38778_o;
  wire [11:0] n38779_o;
  wire [11:0] n38782_o;
  wire [11:0] n38783_o;
  wire [1:0] n38799_o;
  wire n38801_o;
  wire n38803_o;
  wire n38804_o;
  wire [2:0] n38805_o;
  wire [12:0] n38817_o;
  wire [12:0] n38818_o;
  wire [12:0] n38819_o;
  wire [9:0] n38821_o;
  wire [12:0] n38825_o;
  wire [12:0] n38826_o;
  wire [12:0] n38828_o;
  wire [9:0] n38830_o;
  wire [12:0] n38834_o;
  wire [12:0] n38835_o;
  wire n38837_o;
  wire [1:0] n38838_o;
  wire n38840_o;
  wire n38841_o;
  wire [11:0] n38842_o;
  wire [8:0] n38843_o;
  wire [8:0] n38844_o;
  wire [2:0] n38845_o;
  wire [2:0] n38846_o;
  wire [2:0] n38847_o;
  wire n38849_o;
  wire [1:0] n38850_o;
  wire n38852_o;
  wire n38853_o;
  wire n38855_o;
  wire n38856_o;
  wire n38858_o;
  wire [4:0] n38859_o;
  wire [8:0] n38860_o;
  wire [4:0] n38861_o;
  wire [5:0] n38863_o;
  wire [2:0] n38864_o;
  wire [8:0] n38865_o;
  wire [8:0] n38866_o;
  wire [2:0] n38867_o;
  wire [12:0] n38868_o;
  wire n38869_o;
  wire [11:0] n38870_o;
  wire [8:0] n38871_o;
  wire [8:0] n38872_o;
  wire [2:0] n38873_o;
  wire n38875_o;
  wire [4:0] n38876_o;
  wire [8:0] n38877_o;
  wire [4:0] n38878_o;
  wire [5:0] n38880_o;
  wire [2:0] n38881_o;
  wire [8:0] n38882_o;
  wire [8:0] n38883_o;
  wire [2:0] n38884_o;
  wire [11:0] n38885_o;
  wire [11:0] n38886_o;
  wire [11:0] n38887_o;
  wire [11:0] n38888_o;
  wire [11:0] n38889_o;
  wire [11:0] n38892_o;
  wire [11:0] n38893_o;
  wire [1:0] n38909_o;
  wire n38911_o;
  wire n38913_o;
  wire n38914_o;
  wire [2:0] n38915_o;
  wire [12:0] n38927_o;
  wire [12:0] n38928_o;
  wire [12:0] n38929_o;
  wire [9:0] n38931_o;
  wire [12:0] n38935_o;
  wire [12:0] n38936_o;
  wire [12:0] n38938_o;
  wire [9:0] n38940_o;
  wire [12:0] n38944_o;
  wire [12:0] n38945_o;
  wire n38947_o;
  wire [1:0] n38948_o;
  wire n38950_o;
  wire n38951_o;
  wire [11:0] n38952_o;
  wire [8:0] n38953_o;
  wire [8:0] n38954_o;
  wire [2:0] n38955_o;
  wire [2:0] n38956_o;
  wire [2:0] n38957_o;
  wire n38959_o;
  wire [1:0] n38960_o;
  wire n38962_o;
  wire n38963_o;
  wire n38965_o;
  wire n38966_o;
  wire n38968_o;
  wire [4:0] n38969_o;
  wire [8:0] n38970_o;
  wire [4:0] n38971_o;
  wire [5:0] n38973_o;
  wire [2:0] n38974_o;
  wire [8:0] n38975_o;
  wire [8:0] n38976_o;
  wire [2:0] n38977_o;
  wire [12:0] n38978_o;
  wire n38979_o;
  wire [11:0] n38980_o;
  wire [8:0] n38981_o;
  wire [8:0] n38982_o;
  wire [2:0] n38983_o;
  wire n38985_o;
  wire [4:0] n38986_o;
  wire [8:0] n38987_o;
  wire [4:0] n38988_o;
  wire [5:0] n38990_o;
  wire [2:0] n38991_o;
  wire [8:0] n38992_o;
  wire [8:0] n38993_o;
  wire [2:0] n38994_o;
  wire [11:0] n38995_o;
  wire [11:0] n38996_o;
  wire [11:0] n38997_o;
  wire [11:0] n38998_o;
  wire [11:0] n38999_o;
  wire [11:0] n39002_o;
  wire [11:0] n39003_o;
  wire [1:0] n39019_o;
  wire n39021_o;
  wire n39023_o;
  wire n39024_o;
  wire [2:0] n39025_o;
  wire [12:0] n39037_o;
  wire [12:0] n39038_o;
  wire [12:0] n39039_o;
  wire [9:0] n39041_o;
  wire [12:0] n39045_o;
  wire [12:0] n39046_o;
  wire [12:0] n39048_o;
  wire [9:0] n39050_o;
  wire [12:0] n39054_o;
  wire [12:0] n39055_o;
  wire n39057_o;
  wire [1:0] n39058_o;
  wire n39060_o;
  wire n39061_o;
  wire [11:0] n39062_o;
  wire [8:0] n39063_o;
  wire [8:0] n39064_o;
  wire [2:0] n39065_o;
  wire [2:0] n39066_o;
  wire [2:0] n39067_o;
  wire n39069_o;
  wire [1:0] n39070_o;
  wire n39072_o;
  wire n39073_o;
  wire n39075_o;
  wire n39076_o;
  wire n39078_o;
  wire [4:0] n39079_o;
  wire [8:0] n39080_o;
  wire [4:0] n39081_o;
  wire [5:0] n39083_o;
  wire [2:0] n39084_o;
  wire [8:0] n39085_o;
  wire [8:0] n39086_o;
  wire [2:0] n39087_o;
  wire [12:0] n39088_o;
  wire n39089_o;
  wire [11:0] n39090_o;
  wire [8:0] n39091_o;
  wire [8:0] n39092_o;
  wire [2:0] n39093_o;
  wire n39095_o;
  wire [4:0] n39096_o;
  wire [8:0] n39097_o;
  wire [4:0] n39098_o;
  wire [5:0] n39100_o;
  wire [2:0] n39101_o;
  wire [8:0] n39102_o;
  wire [8:0] n39103_o;
  wire [2:0] n39104_o;
  wire [11:0] n39105_o;
  wire [11:0] n39106_o;
  wire [11:0] n39107_o;
  wire [11:0] n39108_o;
  wire [11:0] n39109_o;
  wire [11:0] n39112_o;
  wire [11:0] n39113_o;
  wire n39120_o;
  wire [11:0] n39122_o;
  wire [6:0] n39123_o;
  wire [7:0] n39124_o;
  wire [3:0] n39126_o;
  wire [7:0] n39127_o;
  wire [6:0] n39128_o;
  wire [7:0] n39129_o;
  wire [7:0] n39130_o;
  wire n39133_o;
  wire n39135_o;
  wire n39137_o;
  wire n39139_o;
  wire n39141_o;
  wire [4:0] n39143_o;
  wire [7:0] n39148_o;
  wire [7:0] n39150_o;
  wire [7:0] n39152_o;
  wire [7:0] n39154_o;
  reg [3:0] n39225_q;
  reg [3:0] n39226_q;
  reg [3:0] n39227_q;
  reg [3:0] n39228_q;
  reg [3:0] n39229_q;
  reg [3:0] n39230_q;
  reg n39232_q;
  reg n39233_q;
  reg [12:0] n39234_q;
  reg [12:0] n39235_q;
  reg [12:0] n39236_q;
  reg n39237_q;
  reg n39238_q;
  reg n39239_q;
  reg n39240_q;
  reg n39242_q;
  reg n39243_q;
  reg n39244_q;
  reg n39245_q;
  reg n39246_q;
  reg n39247_q;
  reg [11:0] n39248_q;
  reg n39249_q;
  reg n39250_q;
  reg n39251_q;
  reg [4:0] n39252_q;
  wire [11:0] n39253_o;
  reg [11:0] n39254_q;
  wire [11:0] n39255_o;
  reg [11:0] n39256_q;
  wire [11:0] n39257_o;
  reg [11:0] n39258_q;
  reg n39259_q;
  reg n39260_q;
  reg n39261_q;
  reg n39262_q;
  reg n39263_q;
  reg n39264_q;
  reg [4:0] n39266_q;
  reg [3:0] n39267_q;
  reg [3:0] n39268_q;
  reg [3:0] n39269_q;
  reg [12:0] n39270_q;
  reg [4:0] n39271_q;
  reg [3:0] n39272_q;
  reg [3:0] n39273_q;
  reg [3:0] n39274_q;
  reg [3:0] n39275_q;
  reg [3:0] n39276_q;
  reg [12:0] n39277_q;
  reg [12:0] n39278_q;
  reg [2:0] n39279_q;
  reg [2:0] n39280_q;
  reg [2:0] n39281_q;
  reg [2:0] n39282_q;
  reg n39284_q;
  reg n39285_q;
  reg n39286_q;
  reg n39287_q;
  reg [4:0] n39289_q;
  reg [103:0] n39290_q;
  reg [12:0] n39291_q;
  reg [12:0] n39292_q;
  reg [12:0] n39293_q;
  reg [12:0] n39294_q;
  reg [12:0] n39295_q;
  reg [12:0] n39296_q;
  reg [7:0] n39297_q;
  reg [7:0] n39298_q;
  reg [7:0] n39299_q;
  reg [7:0] n39300_q;
  reg [7:0] n39301_q;
  reg [7:0] n39302_q;
  reg [7:0] n39303_q;
  reg [7:0] n39304_q;
  reg [7:0] n39305_q;
  reg [12:0] n39306_q;
  wire [12:0] n39307_o;
  wire [12:0] n39308_o;
  wire [12:0] n39309_o;
  wire [12:0] n39310_o;
  wire [1:0] n39311_o;
  reg [12:0] n39312_o;
  wire [12:0] n39313_o;
  wire [12:0] n39314_o;
  wire [12:0] n39315_o;
  wire [12:0] n39316_o;
  wire [1:0] n39317_o;
  reg [12:0] n39318_o;
  wire [12:0] n39319_o;
  wire [12:0] n39320_o;
  wire [12:0] n39321_o;
  wire [12:0] n39322_o;
  wire [1:0] n39323_o;
  reg [12:0] n39324_o;
  wire [12:0] n39325_o;
  wire [12:0] n39326_o;
  wire [12:0] n39327_o;
  wire [12:0] n39328_o;
  wire [1:0] n39329_o;
  reg [12:0] n39330_o;
  wire [12:0] n39331_o;
  wire [12:0] n39332_o;
  wire [12:0] n39333_o;
  wire [12:0] n39334_o;
  wire [1:0] n39335_o;
  reg [12:0] n39336_o;
  wire [12:0] n39337_o;
  wire [12:0] n39338_o;
  wire [12:0] n39339_o;
  wire [12:0] n39340_o;
  wire [1:0] n39341_o;
  reg [12:0] n39342_o;
  wire [12:0] n39343_o;
  wire [12:0] n39344_o;
  wire [12:0] n39345_o;
  wire [12:0] n39346_o;
  wire [1:0] n39347_o;
  reg [12:0] n39348_o;
  wire [12:0] n39349_o;
  wire [12:0] n39350_o;
  wire [12:0] n39351_o;
  wire [12:0] n39352_o;
  wire [1:0] n39353_o;
  reg [12:0] n39354_o;
  wire [12:0] n39355_o;
  wire [12:0] n39356_o;
  wire [12:0] n39357_o;
  wire [12:0] n39358_o;
  wire [12:0] n39359_o;
  wire [12:0] n39360_o;
  wire [12:0] n39361_o;
  wire [12:0] n39362_o;
  wire [1:0] n39363_o;
  reg [12:0] n39364_o;
  wire [1:0] n39365_o;
  reg [12:0] n39366_o;
  wire n39367_o;
  wire [12:0] n39368_o;
  wire [12:0] n39369_o;
  wire [12:0] n39370_o;
  wire [12:0] n39371_o;
  wire [12:0] n39372_o;
  wire [12:0] n39373_o;
  wire [12:0] n39374_o;
  wire [12:0] n39375_o;
  wire [12:0] n39376_o;
  wire [1:0] n39377_o;
  reg [12:0] n39378_o;
  wire [1:0] n39379_o;
  reg [12:0] n39380_o;
  wire n39381_o;
  wire [12:0] n39382_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n38441_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n38298_o;
  assign i_x2_out = n38335_o;
  assign result_waddr_out = n38336_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n39225_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n39226_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n39227_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n39228_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n39229_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n39230_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n39232_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n39233_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n39234_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n39235_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n39236_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n39237_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n39238_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n39239_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n39240_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n38339_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n39242_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n39243_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n38337_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n39244_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n38359_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n39245_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n38367_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n39246_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n38372_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n39247_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n39248_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n38341_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n38342_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n38343_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n38344_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n38345_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n38346_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n38347_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n38348_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n38349_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n38350_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n38351_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n38352_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n39249_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n39250_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n39251_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n39252_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n39254_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n39256_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n39258_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n38783_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n38893_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n39003_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n39113_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n39259_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n39260_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n39261_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n39262_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n39263_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n39264_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n38494_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n38495_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n38496_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n38497_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n38498_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n39266_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n39267_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n39268_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n39269_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n39270_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n39271_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n39272_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n39273_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n39274_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n39275_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n39276_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n39277_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n39278_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n39279_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n39280_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n39281_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n39282_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n39284_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n39285_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n39286_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n39287_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n39289_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n39290_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n38374_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n38375_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n39291_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n39292_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n39293_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n39294_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n39295_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n39296_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n38384_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n38394_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n38404_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n39330_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n39336_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n39342_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n38439_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n38431_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n39354_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n39297_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n39298_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n39299_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n39300_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n39301_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n39302_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n39303_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n39304_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n39305_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n39306_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n38269_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n38271_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n38274_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n38276_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n38278_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n38280_o = imu_x1_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38281_o = {n38280_o, n38278_o, n38276_o, n38274_o, n38271_o, n38269_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38283_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38285_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38286_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38287_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n38281_o)
      6'b100000: n38288_o = n38286_o;
      6'b010000: n38288_o = n38285_o;
      6'b001000: n38288_o = 4'b0011;
      6'b000100: n38288_o = instruction_tid_rrr;
      6'b000010: n38288_o = n38283_o;
      6'b000001: n38288_o = 4'b0000;
      default: n38288_o = n38287_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38290_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38292_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38293_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38294_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n38281_o)
      6'b100000: n38295_o = n38293_o;
      6'b010000: n38295_o = n38292_o;
      6'b001000: n38295_o = 9'b000000000;
      6'b000100: n38295_o = 9'b000000000;
      6'b000010: n38295_o = n38290_o;
      6'b000001: n38295_o = 9'b000000000;
      default: n38295_o = n38294_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38298_o = {n38295_o, n38288_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n38306_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n38308_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n38311_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n38313_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n38315_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n38317_o = imu_x2_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38318_o = {n38317_o, n38315_o, n38313_o, n38311_o, n38308_o, n38306_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38320_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38322_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38323_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n38324_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n38318_o)
      6'b100000: n38325_o = n38323_o;
      6'b010000: n38325_o = n38322_o;
      6'b001000: n38325_o = 4'b0011;
      6'b000100: n38325_o = instruction_tid_rrr;
      6'b000010: n38325_o = n38320_o;
      6'b000001: n38325_o = 4'b0000;
      default: n38325_o = n38324_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38327_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38329_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38330_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38331_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n38318_o)
      6'b100000: n38332_o = n38330_o;
      6'b010000: n38332_o = n38329_o;
      6'b001000: n38332_o = 9'b000000000;
      6'b000100: n38332_o = 9'b000000000;
      6'b000010: n38332_o = n38327_o;
      6'b000001: n38332_o = 9'b000000000;
      default: n38332_o = n38331_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n38335_o = {n38332_o, n38325_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n38336_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n38337_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n38338_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n38339_o = instruction_mu_valid_in ? n38338_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n38341_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n38342_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n38343_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n38344_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n38345_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n38346_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n38347_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n38348_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n38349_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n38350_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n38351_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n38352_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n38355_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n38356_o = n38355_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n38357_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n38358_o = n38357_o & n38356_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n38359_o = n38358_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n38363_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n38364_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n38365_o = n38364_o & n38363_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n38366_o = n38365_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n38367_o = n38366_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n38371_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n38372_o = n38371_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n38374_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n38375_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n38376_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n38380_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n38381_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n38382_o = ~n38381_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n38383_o = n38380_o | n38382_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n38384_o = n38383_o ? n39312_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n38386_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n38390_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n38391_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n38392_o = ~n38391_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n38393_o = n38390_o | n38392_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n38394_o = n38393_o ? n39318_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n38396_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n38400_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n38401_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n38402_o = ~n38401_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n38403_o = n38400_o | n38402_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n38404_o = n38403_o ? n39324_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n38406_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n38410_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n38415_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n38423_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n38427_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n38428_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n38429_o = ~n38428_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n38430_o = n38427_o | n38429_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n38431_o = n38430_o ? n39348_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n38433_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n38437_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n38438_o = ~n38437_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n38439_o = n38438_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n38440_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n38441_o = n38440_o ? mu_lane_rrrrrr : n38442_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n38442_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n38445_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n38447_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n38448_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n38449_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n38450_o = ~n38449_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n38451_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n38452_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n38453_o = n38450_o ? n38451_o : n38452_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n38454_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n38455_o = ~n38454_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n38456_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n38457_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n38458_o = n38455_o ? n38456_o : n38457_o;
  assign n38469_o = {n38447_o, n38453_o, n38458_o, n38448_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n38494_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n38495_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n38496_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n38497_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n38498_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n38502_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n38504_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n38508_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n38513_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n38514_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n38516_o = n38514_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n38517_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n38519_o = n38516_o ? n38517_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n38522_o = n38516_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n38524_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n38527_o = n38524_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n38529_o = n38513_o ? n38527_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n38531_o = n38513_o ? n38519_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n38533_o = n38513_o ? n38522_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n38535_o = got_imu_rr ? n38529_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n38537_o = got_imu_rr ? n38531_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n38539_o = got_imu_rr ? n38533_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n38541_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n38689_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n38691_o = n38689_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n38693_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n38694_o = n38691_o | n38693_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n38695_o = mu_x1_parm1[2:0];
  assign n38707_o = {1'b0, mu_x1_parm1};
  assign n38708_o = {10'b0000000000, n38695_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n38709_o = n38694_o ? n38708_o : n38707_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n38711_o = mu_x1_i1_1[9:0];
  assign n38715_o = {n38711_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n38716_o = mu_x1_vector ? n38715_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n38718_o = mu_x1_i0_1 + n38709_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n38720_o = n38718_o[9:0];
  assign n38724_o = {n38720_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n38725_o = mu_x1_vector ? n38724_o : n38718_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n38727_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n38728_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n38730_o = n38728_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n38731_o = n38727_o | n38730_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n38732_o = n38725_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n38733_o = n38732_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n38734_o = ~n38733_o;
  assign n38735_o = n38724_o[2:0];
  assign n38736_o = n38718_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n38737_o = mu_x1_vector ? n38735_o : n38736_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n38739_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n38740_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n38742_o = n38740_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n38743_o = n38739_o | n38742_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n38745_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n38746_o = n38743_o | n38745_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n38748_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n38749_o = n38725_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n38750_o = {n38749_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n38751_o = n38725_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n38753_o = {1'b0, n38751_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n38754_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n38755_o = {n38753_o, n38754_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n38756_o = n38748_o ? n38750_o : n38755_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n38757_o = n38725_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n38758_o = n38716_o + n38725_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n38759_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n38760_o = n38758_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n38761_o = n38760_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n38762_o = ~n38761_o;
  assign n38763_o = n38758_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n38765_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n38766_o = n38758_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n38767_o = {n38766_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n38768_o = n38758_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n38770_o = {1'b0, n38768_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n38771_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n38772_o = {n38770_o, n38771_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n38773_o = n38765_o ? n38767_o : n38772_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n38774_o = n38758_o[2:0];
  assign n38775_o = {n38773_o, n38774_o};
  assign n38776_o = {n38762_o, n38763_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n38777_o = n38759_o ? n38776_o : n38775_o;
  assign n38778_o = {n38756_o, n38757_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n38779_o = n38746_o ? n38778_o : n38777_o;
  assign n38782_o = {n38734_o, n38737_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n38783_o = n38731_o ? n38782_o : n38779_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n38799_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n38801_o = n38799_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n38803_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n38804_o = n38801_o | n38803_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n38805_o = mu_x2_parm1[2:0];
  assign n38817_o = {1'b0, mu_x2_parm1};
  assign n38818_o = {10'b0000000000, n38805_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n38819_o = n38804_o ? n38818_o : n38817_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n38821_o = mu_x2_i1_1[9:0];
  assign n38825_o = {n38821_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n38826_o = mu_x2_vector ? n38825_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n38828_o = mu_x2_i0_1 + n38819_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n38830_o = n38828_o[9:0];
  assign n38834_o = {n38830_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n38835_o = mu_x2_vector ? n38834_o : n38828_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n38837_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n38838_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n38840_o = n38838_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n38841_o = n38837_o | n38840_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n38842_o = n38835_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n38843_o = n38842_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n38844_o = ~n38843_o;
  assign n38845_o = n38834_o[2:0];
  assign n38846_o = n38828_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n38847_o = mu_x2_vector ? n38845_o : n38846_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n38849_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n38850_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n38852_o = n38850_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n38853_o = n38849_o | n38852_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n38855_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n38856_o = n38853_o | n38855_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n38858_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n38859_o = n38835_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n38860_o = {n38859_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n38861_o = n38835_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n38863_o = {1'b0, n38861_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n38864_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n38865_o = {n38863_o, n38864_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n38866_o = n38858_o ? n38860_o : n38865_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n38867_o = n38835_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n38868_o = n38826_o + n38835_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n38869_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n38870_o = n38868_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n38871_o = n38870_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n38872_o = ~n38871_o;
  assign n38873_o = n38868_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n38875_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n38876_o = n38868_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n38877_o = {n38876_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n38878_o = n38868_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n38880_o = {1'b0, n38878_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n38881_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n38882_o = {n38880_o, n38881_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n38883_o = n38875_o ? n38877_o : n38882_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n38884_o = n38868_o[2:0];
  assign n38885_o = {n38883_o, n38884_o};
  assign n38886_o = {n38872_o, n38873_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n38887_o = n38869_o ? n38886_o : n38885_o;
  assign n38888_o = {n38866_o, n38867_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n38889_o = n38856_o ? n38888_o : n38887_o;
  assign n38892_o = {n38844_o, n38847_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n38893_o = n38841_o ? n38892_o : n38889_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n38909_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n38911_o = n38909_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n38913_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n38914_o = n38911_o | n38913_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n38915_o = mu_x3_parm1[2:0];
  assign n38927_o = {1'b0, mu_x3_parm1};
  assign n38928_o = {10'b0000000000, n38915_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n38929_o = n38914_o ? n38928_o : n38927_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n38931_o = mu_x3_i1_1[9:0];
  assign n38935_o = {n38931_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n38936_o = mu_x3_vector ? n38935_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n38938_o = mu_x3_i0_1 + n38929_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n38940_o = n38938_o[9:0];
  assign n38944_o = {n38940_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n38945_o = mu_x3_vector ? n38944_o : n38938_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n38947_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n38948_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n38950_o = n38948_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n38951_o = n38947_o | n38950_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n38952_o = n38945_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n38953_o = n38952_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n38954_o = ~n38953_o;
  assign n38955_o = n38944_o[2:0];
  assign n38956_o = n38938_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n38957_o = mu_x3_vector ? n38955_o : n38956_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n38959_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n38960_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n38962_o = n38960_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n38963_o = n38959_o | n38962_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n38965_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n38966_o = n38963_o | n38965_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n38968_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n38969_o = n38945_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n38970_o = {n38969_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n38971_o = n38945_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n38973_o = {1'b0, n38971_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n38974_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n38975_o = {n38973_o, n38974_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n38976_o = n38968_o ? n38970_o : n38975_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n38977_o = n38945_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n38978_o = n38936_o + n38945_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n38979_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n38980_o = n38978_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n38981_o = n38980_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n38982_o = ~n38981_o;
  assign n38983_o = n38978_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n38985_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n38986_o = n38978_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n38987_o = {n38986_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n38988_o = n38978_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n38990_o = {1'b0, n38988_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n38991_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n38992_o = {n38990_o, n38991_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n38993_o = n38985_o ? n38987_o : n38992_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n38994_o = n38978_o[2:0];
  assign n38995_o = {n38993_o, n38994_o};
  assign n38996_o = {n38982_o, n38983_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n38997_o = n38979_o ? n38996_o : n38995_o;
  assign n38998_o = {n38976_o, n38977_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n38999_o = n38966_o ? n38998_o : n38997_o;
  assign n39002_o = {n38954_o, n38957_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n39003_o = n38951_o ? n39002_o : n38999_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n39019_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n39021_o = n39019_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n39023_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n39024_o = n39021_o | n39023_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n39025_o = mu_y_parm1[2:0];
  assign n39037_o = {1'b0, mu_y_parm1};
  assign n39038_o = {10'b0000000000, n39025_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n39039_o = n39024_o ? n39038_o : n39037_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n39041_o = mu_y_i1_1[9:0];
  assign n39045_o = {n39041_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n39046_o = mu_y_vector ? n39045_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n39048_o = mu_y_i0_1 + n39039_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n39050_o = n39048_o[9:0];
  assign n39054_o = {n39050_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n39055_o = mu_y_vector ? n39054_o : n39048_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n39057_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n39058_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n39060_o = n39058_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n39061_o = n39057_o | n39060_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n39062_o = n39055_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n39063_o = n39062_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n39064_o = ~n39063_o;
  assign n39065_o = n39054_o[2:0];
  assign n39066_o = n39048_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n39067_o = mu_y_vector ? n39065_o : n39066_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n39069_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n39070_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n39072_o = n39070_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n39073_o = n39069_o | n39072_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n39075_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n39076_o = n39073_o | n39075_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n39078_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n39079_o = n39055_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n39080_o = {n39079_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n39081_o = n39055_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n39083_o = {1'b0, n39081_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n39084_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n39085_o = {n39083_o, n39084_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n39086_o = n39078_o ? n39080_o : n39085_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n39087_o = n39055_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n39088_o = n39046_o + n39055_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n39089_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n39090_o = n39088_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n39091_o = n39090_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n39092_o = ~n39091_o;
  assign n39093_o = n39088_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n39095_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n39096_o = n39088_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n39097_o = {n39096_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n39098_o = n39088_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n39100_o = {1'b0, n39098_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n39101_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n39102_o = {n39100_o, n39101_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n39103_o = n39095_o ? n39097_o : n39102_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n39104_o = n39088_o[2:0];
  assign n39105_o = {n39103_o, n39104_o};
  assign n39106_o = {n39092_o, n39093_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n39107_o = n39089_o ? n39106_o : n39105_o;
  assign n39108_o = {n39086_o, n39087_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n39109_o = n39076_o ? n39108_o : n39107_o;
  assign n39112_o = {n39064_o, n39067_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n39113_o = n39061_o ? n39112_o : n39109_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n39120_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n39122_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n39123_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n39124_o = {instruction_vm_in, n39123_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n39126_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n39127_o = {n39126_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n39128_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n39129_o = {instruction_vm_in, n39128_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n39130_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39133_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39135_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39137_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39139_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39141_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39143_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39148_o = instruction_tid_valid_in ? n39130_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39150_o = instruction_tid_valid_in ? n39129_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39152_o = instruction_tid_valid_in ? n39127_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n39154_o = instruction_tid_valid_in ? n39124_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39225_q <= 4'b0000;
    else
      n39225_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39226_q <= 4'b0000;
    else
      n39226_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39227_q <= 4'b0000;
    else
      n39227_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39228_q <= 4'b0000;
    else
      n39228_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39229_q <= 4'b0000;
    else
      n39229_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39230_q <= 4'b0000;
    else
      n39230_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39232_q <= 1'b0;
    else
      n39232_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39233_q <= 1'b0;
    else
      n39233_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39234_q <= 13'b0000000000000;
    else
      n39234_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39235_q <= 13'b0000000000000;
    else
      n39235_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39236_q <= 13'b0000000000000;
    else
      n39236_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39237_q <= 1'b0;
    else
      n39237_q <= n38535_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39238_q <= 1'b0;
    else
      n39238_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39239_q <= 1'b0;
    else
      n39239_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39240_q <= 1'b0;
    else
      n39240_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39242_q <= 1'b0;
    else
      n39242_q <= n39133_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39243_q <= 1'b0;
    else
      n39243_q <= n39135_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39244_q <= 1'b0;
    else
      n39244_q <= n39137_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39245_q <= 1'b0;
    else
      n39245_q <= n39139_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39246_q <= 1'b0;
    else
      n39246_q <= n39141_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39247_q <= 1'b0;
    else
      n39247_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39248_q <= 12'b000000000000;
    else
      n39248_q <= n39122_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39249_q <= 1'b0;
    else
      n39249_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39250_q <= 1'b0;
    else
      n39250_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39251_q <= 1'b0;
    else
      n39251_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39252_q <= 5'b00000;
    else
      n39252_q <= n39143_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n39253_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39254_q <= 12'b000000000000;
    else
      n39254_q <= n39253_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n39255_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39256_q <= 12'b000000000000;
    else
      n39256_q <= n39255_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n39257_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39258_q <= 12'b000000000000;
    else
      n39258_q <= n39257_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39259_q <= 1'b0;
    else
      n39259_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39260_q <= 1'b0;
    else
      n39260_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39261_q <= 1'b0;
    else
      n39261_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39262_q <= 1'b0;
    else
      n39262_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39263_q <= 1'b0;
    else
      n39263_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39264_q <= 1'b0;
    else
      n39264_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39266_q <= 5'b00000;
    else
      n39266_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39267_q <= 4'b0000;
    else
      n39267_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39268_q <= 4'b0000;
    else
      n39268_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39269_q <= 4'b0000;
    else
      n39269_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39270_q <= 13'b0000000000000;
    else
      n39270_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39271_q <= 5'b00000;
    else
      n39271_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39272_q <= 4'b0000;
    else
      n39272_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39273_q <= 4'b0000;
    else
      n39273_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39274_q <= 4'b0000;
    else
      n39274_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39275_q <= 4'b0000;
    else
      n39275_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39276_q <= 4'b0000;
    else
      n39276_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39277_q <= 13'b0000000000000;
    else
      n39277_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39278_q <= 13'b0000000000000;
    else
      n39278_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39279_q <= 3'b000;
    else
      n39279_q <= n38537_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39280_q <= 3'b000;
    else
      n39280_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39281_q <= 3'b000;
    else
      n39281_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39282_q <= 3'b000;
    else
      n39282_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39284_q <= 1'b0;
    else
      n39284_q <= n38539_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39285_q <= 1'b0;
    else
      n39285_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39286_q <= 1'b0;
    else
      n39286_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39287_q <= 1'b0;
    else
      n39287_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39289_q <= 5'b00000;
    else
      n39289_q <= n38541_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n38445_o)
    if (n38445_o)
      n39290_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n39290_q <= n38469_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39291_q <= 13'b0000000000000;
    else
      n39291_q <= n39368_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39292_q <= 13'b0000000000000;
    else
      n39292_q <= n39382_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39293_q <= 13'b0000000000000;
    else
      n39293_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39294_q <= 13'b0000000000000;
    else
      n39294_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39295_q <= 13'b0000000000000;
    else
      n39295_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39296_q <= 13'b0000000000000;
    else
      n39296_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39297_q <= 8'b00000000;
    else
      n39297_q <= n39148_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39298_q <= 8'b00000000;
    else
      n39298_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39299_q <= 8'b00000000;
    else
      n39299_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39300_q <= 8'b00000000;
    else
      n39300_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39301_q <= 8'b00000000;
    else
      n39301_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39302_q <= 8'b00000000;
    else
      n39302_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39303_q <= 8'b00000000;
    else
      n39303_q <= n39150_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39304_q <= 8'b00000000;
    else
      n39304_q <= n39152_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n39120_o)
    if (n39120_o)
      n39305_q <= 8'b00000000;
    else
      n39305_q <= n39154_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n38502_o)
    if (n38502_o)
      n39306_q <= 13'b0000000000000;
    else
      n39306_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n39307_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n39308_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n39309_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n39310_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n39311_o = n38376_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n39311_o)
      2'b00: n39312_o = n39307_o;
      2'b01: n39312_o = n39308_o;
      2'b10: n39312_o = n39309_o;
      2'b11: n39312_o = n39310_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n39313_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n39314_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n39315_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n39316_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n39317_o = n38386_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n39317_o)
      2'b00: n39318_o = n39313_o;
      2'b01: n39318_o = n39314_o;
      2'b10: n39318_o = n39315_o;
      2'b11: n39318_o = n39316_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n39319_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n39320_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n39321_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n39322_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n39323_o = n38396_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n39323_o)
      2'b00: n39324_o = n39319_o;
      2'b01: n39324_o = n39320_o;
      2'b10: n39324_o = n39321_o;
      2'b11: n39324_o = n39322_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n39325_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n39326_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n39327_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n39328_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n39329_o = n38406_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n39329_o)
      2'b00: n39330_o = n39325_o;
      2'b01: n39330_o = n39326_o;
      2'b10: n39330_o = n39327_o;
      2'b11: n39330_o = n39328_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n39331_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n39332_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n39333_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n39334_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n39335_o = n38410_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n39335_o)
      2'b00: n39336_o = n39331_o;
      2'b01: n39336_o = n39332_o;
      2'b10: n39336_o = n39333_o;
      2'b11: n39336_o = n39334_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n39337_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n39338_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n39339_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n39340_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n39341_o = n38415_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n39341_o)
      2'b00: n39342_o = n39337_o;
      2'b01: n39342_o = n39338_o;
      2'b10: n39342_o = n39339_o;
      2'b11: n39342_o = n39340_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n39343_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n39344_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n39345_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n39346_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n39347_o = n38423_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n39347_o)
      2'b00: n39348_o = n39343_o;
      2'b01: n39348_o = n39344_o;
      2'b10: n39348_o = n39345_o;
      2'b11: n39348_o = n39346_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n39349_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n39350_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n39351_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n39352_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n39353_o = n38433_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n39353_o)
      2'b00: n39354_o = n39349_o;
      2'b01: n39354_o = n39350_o;
      2'b10: n39354_o = n39351_o;
      2'b11: n39354_o = n39352_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n39355_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n39356_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n39357_o = iregisters_r[38:26];
  assign n39358_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n39359_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n39360_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n39361_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n39362_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n39363_o = n38504_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n39363_o)
      2'b00: n39364_o = n39355_o;
      2'b01: n39364_o = n39356_o;
      2'b10: n39364_o = n39357_o;
      2'b11: n39364_o = n39358_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n39365_o = n38504_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n39365_o)
      2'b00: n39366_o = n39359_o;
      2'b01: n39366_o = n39360_o;
      2'b10: n39366_o = n39361_o;
      2'b11: n39366_o = n39362_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n39367_o = n38504_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n39368_o = n39367_o ? n39366_o : n39364_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n39369_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n39370_o = iregisters_r[25:13];
  assign n39371_o = iregisters_r[38:26];
  assign n39372_o = iregisters_r[51:39];
  assign n39373_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n39374_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n39375_o = iregisters_r[90:78];
  assign n39376_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n39377_o = n38508_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n39377_o)
      2'b00: n39378_o = n39369_o;
      2'b01: n39378_o = n39370_o;
      2'b10: n39378_o = n39371_o;
      2'b11: n39378_o = n39372_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n39379_o = n38508_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n39379_o)
      2'b00: n39380_o = n39373_o;
      2'b01: n39380_o = n39374_o;
      2'b10: n39380_o = n39375_o;
      2'b11: n39380_o = n39376_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n39381_o = n38508_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n39382_o = n39381_o ? n39380_o : n39378_o;
endmodule

module instr_decoder2_0_2
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n37118_o;
  wire n37120_o;
  wire n37123_o;
  wire n37125_o;
  wire n37127_o;
  wire n37129_o;
  wire [5:0] n37130_o;
  wire [3:0] n37132_o;
  wire [3:0] n37134_o;
  wire [3:0] n37135_o;
  wire [3:0] n37136_o;
  reg [3:0] n37137_o;
  wire [8:0] n37139_o;
  wire [8:0] n37141_o;
  wire [8:0] n37142_o;
  wire [8:0] n37143_o;
  reg [8:0] n37144_o;
  wire [12:0] n37147_o;
  wire n37155_o;
  wire n37157_o;
  wire n37160_o;
  wire n37162_o;
  wire n37164_o;
  wire n37166_o;
  wire [5:0] n37167_o;
  wire [3:0] n37169_o;
  wire [3:0] n37171_o;
  wire [3:0] n37172_o;
  wire [3:0] n37173_o;
  reg [3:0] n37174_o;
  wire [8:0] n37176_o;
  wire [8:0] n37178_o;
  wire [8:0] n37179_o;
  wire [8:0] n37180_o;
  reg [8:0] n37181_o;
  wire [12:0] n37184_o;
  wire [7:0] n37185_o;
  wire n37186_o;
  wire [4:0] n37187_o;
  wire [4:0] n37188_o;
  wire [11:0] n37190_o;
  wire [11:0] n37191_o;
  wire [11:0] n37192_o;
  wire [11:0] n37193_o;
  wire [3:0] n37194_o;
  wire [3:0] n37195_o;
  wire [3:0] n37196_o;
  wire [3:0] n37197_o;
  wire n37198_o;
  wire n37199_o;
  wire n37200_o;
  wire n37201_o;
  wire n37204_o;
  wire n37205_o;
  wire n37206_o;
  wire n37207_o;
  wire n37208_o;
  wire n37212_o;
  wire n37213_o;
  wire n37214_o;
  wire n37215_o;
  wire n37216_o;
  wire n37220_o;
  wire n37221_o;
  wire [51:0] n37223_o;
  wire [51:0] n37224_o;
  wire [1:0] n37225_o;
  wire n37229_o;
  wire n37230_o;
  wire n37231_o;
  wire n37232_o;
  wire [12:0] n37233_o;
  wire [1:0] n37235_o;
  wire n37239_o;
  wire n37240_o;
  wire n37241_o;
  wire n37242_o;
  wire [12:0] n37243_o;
  wire [1:0] n37245_o;
  wire n37249_o;
  wire n37250_o;
  wire n37251_o;
  wire n37252_o;
  wire [12:0] n37253_o;
  wire [1:0] n37255_o;
  wire [1:0] n37259_o;
  wire [1:0] n37264_o;
  wire [1:0] n37272_o;
  wire n37276_o;
  wire n37277_o;
  wire n37278_o;
  wire n37279_o;
  wire [12:0] n37280_o;
  wire [1:0] n37282_o;
  wire n37286_o;
  wire n37287_o;
  wire [12:0] n37288_o;
  wire n37289_o;
  wire [7:0] n37290_o;
  wire [7:0] n37291_o;
  wire n37294_o;
  wire [51:0] n37296_o;
  wire [25:0] n37297_o;
  wire n37298_o;
  wire n37299_o;
  wire [12:0] n37300_o;
  wire [12:0] n37301_o;
  wire [12:0] n37302_o;
  wire n37303_o;
  wire n37304_o;
  wire [12:0] n37305_o;
  wire [12:0] n37306_o;
  wire [12:0] n37307_o;
  wire [103:0] n37318_o;
  wire [4:0] n37343_o;
  wire [3:0] n37344_o;
  wire [3:0] n37345_o;
  wire [3:0] n37346_o;
  wire [12:0] n37347_o;
  wire n37351_o;
  wire [2:0] n37353_o;
  wire [2:0] n37357_o;
  wire n37362_o;
  wire n37363_o;
  wire n37365_o;
  wire [2:0] n37366_o;
  wire [2:0] n37368_o;
  wire n37371_o;
  wire n37373_o;
  wire n37376_o;
  wire n37378_o;
  wire [2:0] n37380_o;
  wire n37382_o;
  wire n37384_o;
  wire [2:0] n37386_o;
  wire n37388_o;
  wire [4:0] n37390_o;
  wire [1:0] n37538_o;
  wire n37540_o;
  wire n37542_o;
  wire n37543_o;
  wire [2:0] n37544_o;
  wire [12:0] n37556_o;
  wire [12:0] n37557_o;
  wire [12:0] n37558_o;
  wire [9:0] n37560_o;
  wire [12:0] n37564_o;
  wire [12:0] n37565_o;
  wire [12:0] n37567_o;
  wire [9:0] n37569_o;
  wire [12:0] n37573_o;
  wire [12:0] n37574_o;
  wire n37576_o;
  wire [1:0] n37577_o;
  wire n37579_o;
  wire n37580_o;
  wire [11:0] n37581_o;
  wire [8:0] n37582_o;
  wire [8:0] n37583_o;
  wire [2:0] n37584_o;
  wire [2:0] n37585_o;
  wire [2:0] n37586_o;
  wire n37588_o;
  wire [1:0] n37589_o;
  wire n37591_o;
  wire n37592_o;
  wire n37594_o;
  wire n37595_o;
  wire n37597_o;
  wire [4:0] n37598_o;
  wire [8:0] n37599_o;
  wire [4:0] n37600_o;
  wire [5:0] n37602_o;
  wire [2:0] n37603_o;
  wire [8:0] n37604_o;
  wire [8:0] n37605_o;
  wire [2:0] n37606_o;
  wire [12:0] n37607_o;
  wire n37608_o;
  wire [11:0] n37609_o;
  wire [8:0] n37610_o;
  wire [8:0] n37611_o;
  wire [2:0] n37612_o;
  wire n37614_o;
  wire [4:0] n37615_o;
  wire [8:0] n37616_o;
  wire [4:0] n37617_o;
  wire [5:0] n37619_o;
  wire [2:0] n37620_o;
  wire [8:0] n37621_o;
  wire [8:0] n37622_o;
  wire [2:0] n37623_o;
  wire [11:0] n37624_o;
  wire [11:0] n37625_o;
  wire [11:0] n37626_o;
  wire [11:0] n37627_o;
  wire [11:0] n37628_o;
  wire [11:0] n37631_o;
  wire [11:0] n37632_o;
  wire [1:0] n37648_o;
  wire n37650_o;
  wire n37652_o;
  wire n37653_o;
  wire [2:0] n37654_o;
  wire [12:0] n37666_o;
  wire [12:0] n37667_o;
  wire [12:0] n37668_o;
  wire [9:0] n37670_o;
  wire [12:0] n37674_o;
  wire [12:0] n37675_o;
  wire [12:0] n37677_o;
  wire [9:0] n37679_o;
  wire [12:0] n37683_o;
  wire [12:0] n37684_o;
  wire n37686_o;
  wire [1:0] n37687_o;
  wire n37689_o;
  wire n37690_o;
  wire [11:0] n37691_o;
  wire [8:0] n37692_o;
  wire [8:0] n37693_o;
  wire [2:0] n37694_o;
  wire [2:0] n37695_o;
  wire [2:0] n37696_o;
  wire n37698_o;
  wire [1:0] n37699_o;
  wire n37701_o;
  wire n37702_o;
  wire n37704_o;
  wire n37705_o;
  wire n37707_o;
  wire [4:0] n37708_o;
  wire [8:0] n37709_o;
  wire [4:0] n37710_o;
  wire [5:0] n37712_o;
  wire [2:0] n37713_o;
  wire [8:0] n37714_o;
  wire [8:0] n37715_o;
  wire [2:0] n37716_o;
  wire [12:0] n37717_o;
  wire n37718_o;
  wire [11:0] n37719_o;
  wire [8:0] n37720_o;
  wire [8:0] n37721_o;
  wire [2:0] n37722_o;
  wire n37724_o;
  wire [4:0] n37725_o;
  wire [8:0] n37726_o;
  wire [4:0] n37727_o;
  wire [5:0] n37729_o;
  wire [2:0] n37730_o;
  wire [8:0] n37731_o;
  wire [8:0] n37732_o;
  wire [2:0] n37733_o;
  wire [11:0] n37734_o;
  wire [11:0] n37735_o;
  wire [11:0] n37736_o;
  wire [11:0] n37737_o;
  wire [11:0] n37738_o;
  wire [11:0] n37741_o;
  wire [11:0] n37742_o;
  wire [1:0] n37758_o;
  wire n37760_o;
  wire n37762_o;
  wire n37763_o;
  wire [2:0] n37764_o;
  wire [12:0] n37776_o;
  wire [12:0] n37777_o;
  wire [12:0] n37778_o;
  wire [9:0] n37780_o;
  wire [12:0] n37784_o;
  wire [12:0] n37785_o;
  wire [12:0] n37787_o;
  wire [9:0] n37789_o;
  wire [12:0] n37793_o;
  wire [12:0] n37794_o;
  wire n37796_o;
  wire [1:0] n37797_o;
  wire n37799_o;
  wire n37800_o;
  wire [11:0] n37801_o;
  wire [8:0] n37802_o;
  wire [8:0] n37803_o;
  wire [2:0] n37804_o;
  wire [2:0] n37805_o;
  wire [2:0] n37806_o;
  wire n37808_o;
  wire [1:0] n37809_o;
  wire n37811_o;
  wire n37812_o;
  wire n37814_o;
  wire n37815_o;
  wire n37817_o;
  wire [4:0] n37818_o;
  wire [8:0] n37819_o;
  wire [4:0] n37820_o;
  wire [5:0] n37822_o;
  wire [2:0] n37823_o;
  wire [8:0] n37824_o;
  wire [8:0] n37825_o;
  wire [2:0] n37826_o;
  wire [12:0] n37827_o;
  wire n37828_o;
  wire [11:0] n37829_o;
  wire [8:0] n37830_o;
  wire [8:0] n37831_o;
  wire [2:0] n37832_o;
  wire n37834_o;
  wire [4:0] n37835_o;
  wire [8:0] n37836_o;
  wire [4:0] n37837_o;
  wire [5:0] n37839_o;
  wire [2:0] n37840_o;
  wire [8:0] n37841_o;
  wire [8:0] n37842_o;
  wire [2:0] n37843_o;
  wire [11:0] n37844_o;
  wire [11:0] n37845_o;
  wire [11:0] n37846_o;
  wire [11:0] n37847_o;
  wire [11:0] n37848_o;
  wire [11:0] n37851_o;
  wire [11:0] n37852_o;
  wire [1:0] n37868_o;
  wire n37870_o;
  wire n37872_o;
  wire n37873_o;
  wire [2:0] n37874_o;
  wire [12:0] n37886_o;
  wire [12:0] n37887_o;
  wire [12:0] n37888_o;
  wire [9:0] n37890_o;
  wire [12:0] n37894_o;
  wire [12:0] n37895_o;
  wire [12:0] n37897_o;
  wire [9:0] n37899_o;
  wire [12:0] n37903_o;
  wire [12:0] n37904_o;
  wire n37906_o;
  wire [1:0] n37907_o;
  wire n37909_o;
  wire n37910_o;
  wire [11:0] n37911_o;
  wire [8:0] n37912_o;
  wire [8:0] n37913_o;
  wire [2:0] n37914_o;
  wire [2:0] n37915_o;
  wire [2:0] n37916_o;
  wire n37918_o;
  wire [1:0] n37919_o;
  wire n37921_o;
  wire n37922_o;
  wire n37924_o;
  wire n37925_o;
  wire n37927_o;
  wire [4:0] n37928_o;
  wire [8:0] n37929_o;
  wire [4:0] n37930_o;
  wire [5:0] n37932_o;
  wire [2:0] n37933_o;
  wire [8:0] n37934_o;
  wire [8:0] n37935_o;
  wire [2:0] n37936_o;
  wire [12:0] n37937_o;
  wire n37938_o;
  wire [11:0] n37939_o;
  wire [8:0] n37940_o;
  wire [8:0] n37941_o;
  wire [2:0] n37942_o;
  wire n37944_o;
  wire [4:0] n37945_o;
  wire [8:0] n37946_o;
  wire [4:0] n37947_o;
  wire [5:0] n37949_o;
  wire [2:0] n37950_o;
  wire [8:0] n37951_o;
  wire [8:0] n37952_o;
  wire [2:0] n37953_o;
  wire [11:0] n37954_o;
  wire [11:0] n37955_o;
  wire [11:0] n37956_o;
  wire [11:0] n37957_o;
  wire [11:0] n37958_o;
  wire [11:0] n37961_o;
  wire [11:0] n37962_o;
  wire n37969_o;
  wire [11:0] n37971_o;
  wire [6:0] n37972_o;
  wire [7:0] n37973_o;
  wire [3:0] n37975_o;
  wire [7:0] n37976_o;
  wire [6:0] n37977_o;
  wire [7:0] n37978_o;
  wire [7:0] n37979_o;
  wire n37982_o;
  wire n37984_o;
  wire n37986_o;
  wire n37988_o;
  wire n37990_o;
  wire [4:0] n37992_o;
  wire [7:0] n37997_o;
  wire [7:0] n37999_o;
  wire [7:0] n38001_o;
  wire [7:0] n38003_o;
  reg [3:0] n38074_q;
  reg [3:0] n38075_q;
  reg [3:0] n38076_q;
  reg [3:0] n38077_q;
  reg [3:0] n38078_q;
  reg [3:0] n38079_q;
  reg n38081_q;
  reg n38082_q;
  reg [12:0] n38083_q;
  reg [12:0] n38084_q;
  reg [12:0] n38085_q;
  reg n38086_q;
  reg n38087_q;
  reg n38088_q;
  reg n38089_q;
  reg n38091_q;
  reg n38092_q;
  reg n38093_q;
  reg n38094_q;
  reg n38095_q;
  reg n38096_q;
  reg [11:0] n38097_q;
  reg n38098_q;
  reg n38099_q;
  reg n38100_q;
  reg [4:0] n38101_q;
  wire [11:0] n38102_o;
  reg [11:0] n38103_q;
  wire [11:0] n38104_o;
  reg [11:0] n38105_q;
  wire [11:0] n38106_o;
  reg [11:0] n38107_q;
  reg n38108_q;
  reg n38109_q;
  reg n38110_q;
  reg n38111_q;
  reg n38112_q;
  reg n38113_q;
  reg [4:0] n38115_q;
  reg [3:0] n38116_q;
  reg [3:0] n38117_q;
  reg [3:0] n38118_q;
  reg [12:0] n38119_q;
  reg [4:0] n38120_q;
  reg [3:0] n38121_q;
  reg [3:0] n38122_q;
  reg [3:0] n38123_q;
  reg [3:0] n38124_q;
  reg [3:0] n38125_q;
  reg [12:0] n38126_q;
  reg [12:0] n38127_q;
  reg [2:0] n38128_q;
  reg [2:0] n38129_q;
  reg [2:0] n38130_q;
  reg [2:0] n38131_q;
  reg n38133_q;
  reg n38134_q;
  reg n38135_q;
  reg n38136_q;
  reg [4:0] n38138_q;
  reg [103:0] n38139_q;
  reg [12:0] n38140_q;
  reg [12:0] n38141_q;
  reg [12:0] n38142_q;
  reg [12:0] n38143_q;
  reg [12:0] n38144_q;
  reg [12:0] n38145_q;
  reg [7:0] n38146_q;
  reg [7:0] n38147_q;
  reg [7:0] n38148_q;
  reg [7:0] n38149_q;
  reg [7:0] n38150_q;
  reg [7:0] n38151_q;
  reg [7:0] n38152_q;
  reg [7:0] n38153_q;
  reg [7:0] n38154_q;
  reg [12:0] n38155_q;
  wire [12:0] n38156_o;
  wire [12:0] n38157_o;
  wire [12:0] n38158_o;
  wire [12:0] n38159_o;
  wire [1:0] n38160_o;
  reg [12:0] n38161_o;
  wire [12:0] n38162_o;
  wire [12:0] n38163_o;
  wire [12:0] n38164_o;
  wire [12:0] n38165_o;
  wire [1:0] n38166_o;
  reg [12:0] n38167_o;
  wire [12:0] n38168_o;
  wire [12:0] n38169_o;
  wire [12:0] n38170_o;
  wire [12:0] n38171_o;
  wire [1:0] n38172_o;
  reg [12:0] n38173_o;
  wire [12:0] n38174_o;
  wire [12:0] n38175_o;
  wire [12:0] n38176_o;
  wire [12:0] n38177_o;
  wire [1:0] n38178_o;
  reg [12:0] n38179_o;
  wire [12:0] n38180_o;
  wire [12:0] n38181_o;
  wire [12:0] n38182_o;
  wire [12:0] n38183_o;
  wire [1:0] n38184_o;
  reg [12:0] n38185_o;
  wire [12:0] n38186_o;
  wire [12:0] n38187_o;
  wire [12:0] n38188_o;
  wire [12:0] n38189_o;
  wire [1:0] n38190_o;
  reg [12:0] n38191_o;
  wire [12:0] n38192_o;
  wire [12:0] n38193_o;
  wire [12:0] n38194_o;
  wire [12:0] n38195_o;
  wire [1:0] n38196_o;
  reg [12:0] n38197_o;
  wire [12:0] n38198_o;
  wire [12:0] n38199_o;
  wire [12:0] n38200_o;
  wire [12:0] n38201_o;
  wire [1:0] n38202_o;
  reg [12:0] n38203_o;
  wire [12:0] n38204_o;
  wire [12:0] n38205_o;
  wire [12:0] n38206_o;
  wire [12:0] n38207_o;
  wire [12:0] n38208_o;
  wire [12:0] n38209_o;
  wire [12:0] n38210_o;
  wire [12:0] n38211_o;
  wire [1:0] n38212_o;
  reg [12:0] n38213_o;
  wire [1:0] n38214_o;
  reg [12:0] n38215_o;
  wire n38216_o;
  wire [12:0] n38217_o;
  wire [12:0] n38218_o;
  wire [12:0] n38219_o;
  wire [12:0] n38220_o;
  wire [12:0] n38221_o;
  wire [12:0] n38222_o;
  wire [12:0] n38223_o;
  wire [12:0] n38224_o;
  wire [12:0] n38225_o;
  wire [1:0] n38226_o;
  reg [12:0] n38227_o;
  wire [1:0] n38228_o;
  reg [12:0] n38229_o;
  wire n38230_o;
  wire [12:0] n38231_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n37290_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n37147_o;
  assign i_x2_out = n37184_o;
  assign result_waddr_out = n37185_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n38074_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n38075_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n38076_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n38077_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n38078_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n38079_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n38081_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n38082_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n38083_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n38084_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n38085_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n38086_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n38087_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n38088_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n38089_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n37188_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n38091_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n38092_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n37186_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n38093_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n37208_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n38094_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n37216_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n38095_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n37221_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n38096_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n38097_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n37190_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n37191_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n37192_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n37193_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n37194_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n37195_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n37196_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n37197_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n37198_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n37199_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n37200_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n37201_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n38098_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n38099_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n38100_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n38101_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n38103_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n38105_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n38107_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n37632_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n37742_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n37852_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n37962_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n38108_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n38109_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n38110_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n38111_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n38112_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n38113_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n37343_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n37344_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n37345_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n37346_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n37347_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n38115_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n38116_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n38117_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n38118_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n38119_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n38120_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n38121_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n38122_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n38123_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n38124_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n38125_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n38126_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n38127_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n38128_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n38129_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n38130_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n38131_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n38133_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n38134_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n38135_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n38136_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n38138_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n38139_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n37223_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n37224_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n38140_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n38141_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n38142_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n38143_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n38144_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n38145_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n37233_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n37243_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n37253_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n38179_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n38185_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n38191_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n37288_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n37280_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n38203_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n38146_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n38147_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n38148_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n38149_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n38150_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n38151_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n38152_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n38153_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n38154_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n38155_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n37118_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n37120_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n37123_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n37125_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n37127_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n37129_o = imu_x1_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37130_o = {n37129_o, n37127_o, n37125_o, n37123_o, n37120_o, n37118_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37132_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37134_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37135_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37136_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n37130_o)
      6'b100000: n37137_o = n37135_o;
      6'b010000: n37137_o = n37134_o;
      6'b001000: n37137_o = 4'b0010;
      6'b000100: n37137_o = instruction_tid_rrr;
      6'b000010: n37137_o = n37132_o;
      6'b000001: n37137_o = 4'b0000;
      default: n37137_o = n37136_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37139_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37141_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37142_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37143_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n37130_o)
      6'b100000: n37144_o = n37142_o;
      6'b010000: n37144_o = n37141_o;
      6'b001000: n37144_o = 9'b000000000;
      6'b000100: n37144_o = 9'b000000000;
      6'b000010: n37144_o = n37139_o;
      6'b000001: n37144_o = 9'b000000000;
      default: n37144_o = n37143_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37147_o = {n37144_o, n37137_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n37155_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n37157_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n37160_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n37162_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n37164_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n37166_o = imu_x2_parm_rrr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37167_o = {n37166_o, n37164_o, n37162_o, n37160_o, n37157_o, n37155_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37169_o = imu_const_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37171_o = result_r[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37172_o = lane_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:1  */
  assign n37173_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n37167_o)
      6'b100000: n37174_o = n37172_o;
      6'b010000: n37174_o = n37171_o;
      6'b001000: n37174_o = 4'b0010;
      6'b000100: n37174_o = instruction_tid_rrr;
      6'b000010: n37174_o = n37169_o;
      6'b000001: n37174_o = 4'b0000;
      default: n37174_o = n37173_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37176_o = imu_const_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37178_o = result_r[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37179_o = lane_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37180_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n37167_o)
      6'b100000: n37181_o = n37179_o;
      6'b010000: n37181_o = n37178_o;
      6'b001000: n37181_o = 9'b000000000;
      6'b000100: n37181_o = 9'b000000000;
      6'b000010: n37181_o = n37176_o;
      6'b000001: n37181_o = 9'b000000000;
      default: n37181_o = n37180_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:5  */
  assign n37184_o = {n37181_o, n37174_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n37185_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n37186_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n37187_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n37188_o = instruction_mu_valid_in ? n37187_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n37190_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n37191_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n37192_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n37193_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n37194_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n37195_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n37196_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n37197_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n37198_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n37199_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n37200_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n37201_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n37204_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n37205_o = n37204_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n37206_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n37207_o = n37206_o & n37205_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n37208_o = n37207_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n37212_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n37213_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n37214_o = n37213_o & n37212_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n37215_o = n37214_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n37216_o = n37215_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n37220_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n37221_o = n37220_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n37223_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n37224_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n37225_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n37229_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n37230_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n37231_o = ~n37230_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n37232_o = n37229_o | n37231_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n37233_o = n37232_o ? n38161_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n37235_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n37239_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n37240_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n37241_o = ~n37240_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n37242_o = n37239_o | n37241_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n37243_o = n37242_o ? n38167_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n37245_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n37249_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n37250_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n37251_o = ~n37250_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n37252_o = n37249_o | n37251_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n37253_o = n37252_o ? n38173_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n37255_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n37259_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n37264_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n37272_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n37276_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n37277_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n37278_o = ~n37277_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n37279_o = n37276_o | n37278_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n37280_o = n37279_o ? n38197_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n37282_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n37286_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n37287_o = ~n37286_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n37288_o = n37287_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n37289_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n37290_o = n37289_o ? mu_lane_rrrrrr : n37291_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n37291_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n37294_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n37296_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n37297_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n37298_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n37299_o = ~n37298_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n37300_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n37301_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n37302_o = n37299_o ? n37300_o : n37301_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n37303_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n37304_o = ~n37303_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n37305_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n37306_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n37307_o = n37304_o ? n37305_o : n37306_o;
  assign n37318_o = {n37296_o, n37302_o, n37307_o, n37297_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n37343_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n37344_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n37345_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n37346_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n37347_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n37351_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n37353_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n37357_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n37362_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n37363_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n37365_o = n37363_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n37366_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n37368_o = n37365_o ? n37366_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n37371_o = n37365_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n37373_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n37376_o = n37373_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n37378_o = n37362_o ? n37376_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n37380_o = n37362_o ? n37368_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n37382_o = n37362_o ? n37371_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n37384_o = got_imu_rr ? n37378_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n37386_o = got_imu_rr ? n37380_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n37388_o = got_imu_rr ? n37382_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n37390_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n37538_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n37540_o = n37538_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n37542_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n37543_o = n37540_o | n37542_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n37544_o = mu_x1_parm1[2:0];
  assign n37556_o = {1'b0, mu_x1_parm1};
  assign n37557_o = {10'b0000000000, n37544_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n37558_o = n37543_o ? n37557_o : n37556_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n37560_o = mu_x1_i1_1[9:0];
  assign n37564_o = {n37560_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n37565_o = mu_x1_vector ? n37564_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n37567_o = mu_x1_i0_1 + n37558_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n37569_o = n37567_o[9:0];
  assign n37573_o = {n37569_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37574_o = mu_x1_vector ? n37573_o : n37567_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n37576_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n37577_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n37579_o = n37577_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n37580_o = n37576_o | n37579_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n37581_o = n37574_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n37582_o = n37581_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n37583_o = ~n37582_o;
  assign n37584_o = n37573_o[2:0];
  assign n37585_o = n37567_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37586_o = mu_x1_vector ? n37584_o : n37585_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n37588_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n37589_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n37591_o = n37589_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n37592_o = n37588_o | n37591_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n37594_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n37595_o = n37592_o | n37594_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n37597_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n37598_o = n37574_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n37599_o = {n37598_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n37600_o = n37574_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n37602_o = {1'b0, n37600_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n37603_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n37604_o = {n37602_o, n37603_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n37605_o = n37597_o ? n37599_o : n37604_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n37606_o = n37574_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n37607_o = n37565_o + n37574_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n37608_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n37609_o = n37607_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n37610_o = n37609_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n37611_o = ~n37610_o;
  assign n37612_o = n37607_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n37614_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n37615_o = n37607_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n37616_o = {n37615_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n37617_o = n37607_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n37619_o = {1'b0, n37617_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n37620_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n37621_o = {n37619_o, n37620_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n37622_o = n37614_o ? n37616_o : n37621_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n37623_o = n37607_o[2:0];
  assign n37624_o = {n37622_o, n37623_o};
  assign n37625_o = {n37611_o, n37612_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n37626_o = n37608_o ? n37625_o : n37624_o;
  assign n37627_o = {n37605_o, n37606_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n37628_o = n37595_o ? n37627_o : n37626_o;
  assign n37631_o = {n37583_o, n37586_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n37632_o = n37580_o ? n37631_o : n37628_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n37648_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n37650_o = n37648_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n37652_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n37653_o = n37650_o | n37652_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n37654_o = mu_x2_parm1[2:0];
  assign n37666_o = {1'b0, mu_x2_parm1};
  assign n37667_o = {10'b0000000000, n37654_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n37668_o = n37653_o ? n37667_o : n37666_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n37670_o = mu_x2_i1_1[9:0];
  assign n37674_o = {n37670_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n37675_o = mu_x2_vector ? n37674_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n37677_o = mu_x2_i0_1 + n37668_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n37679_o = n37677_o[9:0];
  assign n37683_o = {n37679_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37684_o = mu_x2_vector ? n37683_o : n37677_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n37686_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n37687_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n37689_o = n37687_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n37690_o = n37686_o | n37689_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n37691_o = n37684_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n37692_o = n37691_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n37693_o = ~n37692_o;
  assign n37694_o = n37683_o[2:0];
  assign n37695_o = n37677_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37696_o = mu_x2_vector ? n37694_o : n37695_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n37698_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n37699_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n37701_o = n37699_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n37702_o = n37698_o | n37701_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n37704_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n37705_o = n37702_o | n37704_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n37707_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n37708_o = n37684_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n37709_o = {n37708_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n37710_o = n37684_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n37712_o = {1'b0, n37710_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n37713_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n37714_o = {n37712_o, n37713_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n37715_o = n37707_o ? n37709_o : n37714_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n37716_o = n37684_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n37717_o = n37675_o + n37684_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n37718_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n37719_o = n37717_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n37720_o = n37719_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n37721_o = ~n37720_o;
  assign n37722_o = n37717_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n37724_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n37725_o = n37717_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n37726_o = {n37725_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n37727_o = n37717_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n37729_o = {1'b0, n37727_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n37730_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n37731_o = {n37729_o, n37730_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n37732_o = n37724_o ? n37726_o : n37731_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n37733_o = n37717_o[2:0];
  assign n37734_o = {n37732_o, n37733_o};
  assign n37735_o = {n37721_o, n37722_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n37736_o = n37718_o ? n37735_o : n37734_o;
  assign n37737_o = {n37715_o, n37716_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n37738_o = n37705_o ? n37737_o : n37736_o;
  assign n37741_o = {n37693_o, n37696_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n37742_o = n37690_o ? n37741_o : n37738_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n37758_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n37760_o = n37758_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n37762_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n37763_o = n37760_o | n37762_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n37764_o = mu_x3_parm1[2:0];
  assign n37776_o = {1'b0, mu_x3_parm1};
  assign n37777_o = {10'b0000000000, n37764_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n37778_o = n37763_o ? n37777_o : n37776_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n37780_o = mu_x3_i1_1[9:0];
  assign n37784_o = {n37780_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n37785_o = mu_x3_vector ? n37784_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n37787_o = mu_x3_i0_1 + n37778_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n37789_o = n37787_o[9:0];
  assign n37793_o = {n37789_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37794_o = mu_x3_vector ? n37793_o : n37787_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n37796_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n37797_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n37799_o = n37797_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n37800_o = n37796_o | n37799_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n37801_o = n37794_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n37802_o = n37801_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n37803_o = ~n37802_o;
  assign n37804_o = n37793_o[2:0];
  assign n37805_o = n37787_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37806_o = mu_x3_vector ? n37804_o : n37805_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n37808_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n37809_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n37811_o = n37809_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n37812_o = n37808_o | n37811_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n37814_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n37815_o = n37812_o | n37814_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n37817_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n37818_o = n37794_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n37819_o = {n37818_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n37820_o = n37794_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n37822_o = {1'b0, n37820_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n37823_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n37824_o = {n37822_o, n37823_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n37825_o = n37817_o ? n37819_o : n37824_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n37826_o = n37794_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n37827_o = n37785_o + n37794_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n37828_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n37829_o = n37827_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n37830_o = n37829_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n37831_o = ~n37830_o;
  assign n37832_o = n37827_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n37834_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n37835_o = n37827_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n37836_o = {n37835_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n37837_o = n37827_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n37839_o = {1'b0, n37837_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n37840_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n37841_o = {n37839_o, n37840_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n37842_o = n37834_o ? n37836_o : n37841_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n37843_o = n37827_o[2:0];
  assign n37844_o = {n37842_o, n37843_o};
  assign n37845_o = {n37831_o, n37832_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n37846_o = n37828_o ? n37845_o : n37844_o;
  assign n37847_o = {n37825_o, n37826_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n37848_o = n37815_o ? n37847_o : n37846_o;
  assign n37851_o = {n37803_o, n37806_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n37852_o = n37800_o ? n37851_o : n37848_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n37868_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n37870_o = n37868_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n37872_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n37873_o = n37870_o | n37872_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n37874_o = mu_y_parm1[2:0];
  assign n37886_o = {1'b0, mu_y_parm1};
  assign n37887_o = {10'b0000000000, n37874_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n37888_o = n37873_o ? n37887_o : n37886_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n37890_o = mu_y_i1_1[9:0];
  assign n37894_o = {n37890_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n37895_o = mu_y_vector ? n37894_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n37897_o = mu_y_i0_1 + n37888_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n37899_o = n37897_o[9:0];
  assign n37903_o = {n37899_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37904_o = mu_y_vector ? n37903_o : n37897_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n37906_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n37907_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n37909_o = n37907_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n37910_o = n37906_o | n37909_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n37911_o = n37904_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n37912_o = n37911_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n37913_o = ~n37912_o;
  assign n37914_o = n37903_o[2:0];
  assign n37915_o = n37897_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n37916_o = mu_y_vector ? n37914_o : n37915_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n37918_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n37919_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n37921_o = n37919_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n37922_o = n37918_o | n37921_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n37924_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n37925_o = n37922_o | n37924_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n37927_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n37928_o = n37904_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n37929_o = {n37928_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n37930_o = n37904_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n37932_o = {1'b0, n37930_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n37933_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n37934_o = {n37932_o, n37933_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n37935_o = n37927_o ? n37929_o : n37934_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n37936_o = n37904_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n37937_o = n37895_o + n37904_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n37938_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n37939_o = n37937_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n37940_o = n37939_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n37941_o = ~n37940_o;
  assign n37942_o = n37937_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n37944_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n37945_o = n37937_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n37946_o = {n37945_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n37947_o = n37937_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n37949_o = {1'b0, n37947_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n37950_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n37951_o = {n37949_o, n37950_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n37952_o = n37944_o ? n37946_o : n37951_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n37953_o = n37937_o[2:0];
  assign n37954_o = {n37952_o, n37953_o};
  assign n37955_o = {n37941_o, n37942_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n37956_o = n37938_o ? n37955_o : n37954_o;
  assign n37957_o = {n37935_o, n37936_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n37958_o = n37925_o ? n37957_o : n37956_o;
  assign n37961_o = {n37913_o, n37916_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n37962_o = n37910_o ? n37961_o : n37958_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n37969_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n37971_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n37972_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n37973_o = {instruction_vm_in, n37972_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n37975_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n37976_o = {n37975_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n37977_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n37978_o = {instruction_vm_in, n37977_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n37979_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37982_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37984_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37986_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37988_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37990_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37992_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37997_o = instruction_tid_valid_in ? n37979_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n37999_o = instruction_tid_valid_in ? n37978_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n38001_o = instruction_tid_valid_in ? n37976_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n38003_o = instruction_tid_valid_in ? n37973_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38074_q <= 4'b0000;
    else
      n38074_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38075_q <= 4'b0000;
    else
      n38075_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38076_q <= 4'b0000;
    else
      n38076_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38077_q <= 4'b0000;
    else
      n38077_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38078_q <= 4'b0000;
    else
      n38078_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38079_q <= 4'b0000;
    else
      n38079_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38081_q <= 1'b0;
    else
      n38081_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38082_q <= 1'b0;
    else
      n38082_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38083_q <= 13'b0000000000000;
    else
      n38083_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38084_q <= 13'b0000000000000;
    else
      n38084_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38085_q <= 13'b0000000000000;
    else
      n38085_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38086_q <= 1'b0;
    else
      n38086_q <= n37384_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38087_q <= 1'b0;
    else
      n38087_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38088_q <= 1'b0;
    else
      n38088_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38089_q <= 1'b0;
    else
      n38089_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38091_q <= 1'b0;
    else
      n38091_q <= n37982_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38092_q <= 1'b0;
    else
      n38092_q <= n37984_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38093_q <= 1'b0;
    else
      n38093_q <= n37986_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38094_q <= 1'b0;
    else
      n38094_q <= n37988_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38095_q <= 1'b0;
    else
      n38095_q <= n37990_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38096_q <= 1'b0;
    else
      n38096_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38097_q <= 12'b000000000000;
    else
      n38097_q <= n37971_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38098_q <= 1'b0;
    else
      n38098_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38099_q <= 1'b0;
    else
      n38099_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38100_q <= 1'b0;
    else
      n38100_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38101_q <= 5'b00000;
    else
      n38101_q <= n37992_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n38102_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38103_q <= 12'b000000000000;
    else
      n38103_q <= n38102_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n38104_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38105_q <= 12'b000000000000;
    else
      n38105_q <= n38104_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n38106_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38107_q <= 12'b000000000000;
    else
      n38107_q <= n38106_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38108_q <= 1'b0;
    else
      n38108_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38109_q <= 1'b0;
    else
      n38109_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38110_q <= 1'b0;
    else
      n38110_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38111_q <= 1'b0;
    else
      n38111_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38112_q <= 1'b0;
    else
      n38112_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38113_q <= 1'b0;
    else
      n38113_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38115_q <= 5'b00000;
    else
      n38115_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38116_q <= 4'b0000;
    else
      n38116_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38117_q <= 4'b0000;
    else
      n38117_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38118_q <= 4'b0000;
    else
      n38118_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38119_q <= 13'b0000000000000;
    else
      n38119_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38120_q <= 5'b00000;
    else
      n38120_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38121_q <= 4'b0000;
    else
      n38121_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38122_q <= 4'b0000;
    else
      n38122_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38123_q <= 4'b0000;
    else
      n38123_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38124_q <= 4'b0000;
    else
      n38124_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38125_q <= 4'b0000;
    else
      n38125_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38126_q <= 13'b0000000000000;
    else
      n38126_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38127_q <= 13'b0000000000000;
    else
      n38127_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38128_q <= 3'b000;
    else
      n38128_q <= n37386_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38129_q <= 3'b000;
    else
      n38129_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38130_q <= 3'b000;
    else
      n38130_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38131_q <= 3'b000;
    else
      n38131_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38133_q <= 1'b0;
    else
      n38133_q <= n37388_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38134_q <= 1'b0;
    else
      n38134_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38135_q <= 1'b0;
    else
      n38135_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38136_q <= 1'b0;
    else
      n38136_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38138_q <= 5'b00000;
    else
      n38138_q <= n37390_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n37294_o)
    if (n37294_o)
      n38139_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n38139_q <= n37318_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38140_q <= 13'b0000000000000;
    else
      n38140_q <= n38217_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38141_q <= 13'b0000000000000;
    else
      n38141_q <= n38231_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38142_q <= 13'b0000000000000;
    else
      n38142_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38143_q <= 13'b0000000000000;
    else
      n38143_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38144_q <= 13'b0000000000000;
    else
      n38144_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38145_q <= 13'b0000000000000;
    else
      n38145_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38146_q <= 8'b00000000;
    else
      n38146_q <= n37997_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38147_q <= 8'b00000000;
    else
      n38147_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38148_q <= 8'b00000000;
    else
      n38148_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38149_q <= 8'b00000000;
    else
      n38149_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38150_q <= 8'b00000000;
    else
      n38150_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38151_q <= 8'b00000000;
    else
      n38151_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38152_q <= 8'b00000000;
    else
      n38152_q <= n37999_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38153_q <= 8'b00000000;
    else
      n38153_q <= n38001_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n37969_o)
    if (n37969_o)
      n38154_q <= 8'b00000000;
    else
      n38154_q <= n38003_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n37351_o)
    if (n37351_o)
      n38155_q <= 13'b0000000000000;
    else
      n38155_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n38156_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n38157_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n38158_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n38159_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n38160_o = n37225_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n38160_o)
      2'b00: n38161_o = n38156_o;
      2'b01: n38161_o = n38157_o;
      2'b10: n38161_o = n38158_o;
      2'b11: n38161_o = n38159_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n38162_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n38163_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n38164_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n38165_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n38166_o = n37235_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n38166_o)
      2'b00: n38167_o = n38162_o;
      2'b01: n38167_o = n38163_o;
      2'b10: n38167_o = n38164_o;
      2'b11: n38167_o = n38165_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n38168_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n38169_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n38170_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n38171_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n38172_o = n37245_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n38172_o)
      2'b00: n38173_o = n38168_o;
      2'b01: n38173_o = n38169_o;
      2'b10: n38173_o = n38170_o;
      2'b11: n38173_o = n38171_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n38174_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n38175_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n38176_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n38177_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n38178_o = n37255_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n38178_o)
      2'b00: n38179_o = n38174_o;
      2'b01: n38179_o = n38175_o;
      2'b10: n38179_o = n38176_o;
      2'b11: n38179_o = n38177_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n38180_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n38181_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n38182_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n38183_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n38184_o = n37259_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n38184_o)
      2'b00: n38185_o = n38180_o;
      2'b01: n38185_o = n38181_o;
      2'b10: n38185_o = n38182_o;
      2'b11: n38185_o = n38183_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n38186_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n38187_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n38188_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n38189_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n38190_o = n37264_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n38190_o)
      2'b00: n38191_o = n38186_o;
      2'b01: n38191_o = n38187_o;
      2'b10: n38191_o = n38188_o;
      2'b11: n38191_o = n38189_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n38192_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n38193_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n38194_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n38195_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n38196_o = n37272_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n38196_o)
      2'b00: n38197_o = n38192_o;
      2'b01: n38197_o = n38193_o;
      2'b10: n38197_o = n38194_o;
      2'b11: n38197_o = n38195_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n38198_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n38199_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n38200_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n38201_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n38202_o = n37282_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n38202_o)
      2'b00: n38203_o = n38198_o;
      2'b01: n38203_o = n38199_o;
      2'b10: n38203_o = n38200_o;
      2'b11: n38203_o = n38201_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n38204_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n38205_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n38206_o = iregisters_r[38:26];
  assign n38207_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n38208_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n38209_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n38210_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n38211_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n38212_o = n37353_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n38212_o)
      2'b00: n38213_o = n38204_o;
      2'b01: n38213_o = n38205_o;
      2'b10: n38213_o = n38206_o;
      2'b11: n38213_o = n38207_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n38214_o = n37353_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n38214_o)
      2'b00: n38215_o = n38208_o;
      2'b01: n38215_o = n38209_o;
      2'b10: n38215_o = n38210_o;
      2'b11: n38215_o = n38211_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n38216_o = n37353_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n38217_o = n38216_o ? n38215_o : n38213_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n38218_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n38219_o = iregisters_r[25:13];
  assign n38220_o = iregisters_r[38:26];
  assign n38221_o = iregisters_r[51:39];
  assign n38222_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n38223_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n38224_o = iregisters_r[90:78];
  assign n38225_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n38226_o = n37357_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n38226_o)
      2'b00: n38227_o = n38218_o;
      2'b01: n38227_o = n38219_o;
      2'b10: n38227_o = n38220_o;
      2'b11: n38227_o = n38221_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n38228_o = n37357_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n38228_o)
      2'b00: n38229_o = n38222_o;
      2'b01: n38229_o = n38223_o;
      2'b10: n38229_o = n38224_o;
      2'b11: n38229_o = n38225_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n38230_o = n37357_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n38231_o = n38230_o ? n38229_o : n38227_o;
endmodule

module instr_decoder2_0_1
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n35967_o;
  wire n35969_o;
  wire n35972_o;
  wire n35974_o;
  wire n35976_o;
  wire n35978_o;
  wire [5:0] n35979_o;
  wire [3:0] n35981_o;
  wire [3:0] n35983_o;
  wire [3:0] n35984_o;
  wire [3:0] n35985_o;
  reg [3:0] n35986_o;
  wire [8:0] n35988_o;
  wire [8:0] n35990_o;
  wire [8:0] n35991_o;
  wire [8:0] n35992_o;
  reg [8:0] n35993_o;
  wire [12:0] n35996_o;
  wire n36004_o;
  wire n36006_o;
  wire n36009_o;
  wire n36011_o;
  wire n36013_o;
  wire n36015_o;
  wire [5:0] n36016_o;
  wire [3:0] n36018_o;
  wire [3:0] n36020_o;
  wire [3:0] n36021_o;
  wire [3:0] n36022_o;
  reg [3:0] n36023_o;
  wire [8:0] n36025_o;
  wire [8:0] n36027_o;
  wire [8:0] n36028_o;
  wire [8:0] n36029_o;
  reg [8:0] n36030_o;
  wire [12:0] n36033_o;
  wire [7:0] n36034_o;
  wire n36035_o;
  wire [4:0] n36036_o;
  wire [4:0] n36037_o;
  wire [11:0] n36039_o;
  wire [11:0] n36040_o;
  wire [11:0] n36041_o;
  wire [11:0] n36042_o;
  wire [3:0] n36043_o;
  wire [3:0] n36044_o;
  wire [3:0] n36045_o;
  wire [3:0] n36046_o;
  wire n36047_o;
  wire n36048_o;
  wire n36049_o;
  wire n36050_o;
  wire n36053_o;
  wire n36054_o;
  wire n36055_o;
  wire n36056_o;
  wire n36057_o;
  wire n36061_o;
  wire n36062_o;
  wire n36063_o;
  wire n36064_o;
  wire n36065_o;
  wire n36069_o;
  wire n36070_o;
  wire [51:0] n36072_o;
  wire [51:0] n36073_o;
  wire [1:0] n36074_o;
  wire n36078_o;
  wire n36079_o;
  wire n36080_o;
  wire n36081_o;
  wire [12:0] n36082_o;
  wire [1:0] n36084_o;
  wire n36088_o;
  wire n36089_o;
  wire n36090_o;
  wire n36091_o;
  wire [12:0] n36092_o;
  wire [1:0] n36094_o;
  wire n36098_o;
  wire n36099_o;
  wire n36100_o;
  wire n36101_o;
  wire [12:0] n36102_o;
  wire [1:0] n36104_o;
  wire [1:0] n36108_o;
  wire [1:0] n36113_o;
  wire [1:0] n36121_o;
  wire n36125_o;
  wire n36126_o;
  wire n36127_o;
  wire n36128_o;
  wire [12:0] n36129_o;
  wire [1:0] n36131_o;
  wire n36135_o;
  wire n36136_o;
  wire [12:0] n36137_o;
  wire n36138_o;
  wire [7:0] n36139_o;
  wire [7:0] n36140_o;
  wire n36143_o;
  wire [51:0] n36145_o;
  wire [25:0] n36146_o;
  wire n36147_o;
  wire n36148_o;
  wire [12:0] n36149_o;
  wire [12:0] n36150_o;
  wire [12:0] n36151_o;
  wire n36152_o;
  wire n36153_o;
  wire [12:0] n36154_o;
  wire [12:0] n36155_o;
  wire [12:0] n36156_o;
  wire [103:0] n36167_o;
  wire [4:0] n36192_o;
  wire [3:0] n36193_o;
  wire [3:0] n36194_o;
  wire [3:0] n36195_o;
  wire [12:0] n36196_o;
  wire n36200_o;
  wire [2:0] n36202_o;
  wire [2:0] n36206_o;
  wire n36211_o;
  wire n36212_o;
  wire n36214_o;
  wire [2:0] n36215_o;
  wire [2:0] n36217_o;
  wire n36220_o;
  wire n36222_o;
  wire n36225_o;
  wire n36227_o;
  wire [2:0] n36229_o;
  wire n36231_o;
  wire n36233_o;
  wire [2:0] n36235_o;
  wire n36237_o;
  wire [4:0] n36239_o;
  wire [1:0] n36387_o;
  wire n36389_o;
  wire n36391_o;
  wire n36392_o;
  wire [2:0] n36393_o;
  wire [12:0] n36405_o;
  wire [12:0] n36406_o;
  wire [12:0] n36407_o;
  wire [9:0] n36409_o;
  wire [12:0] n36413_o;
  wire [12:0] n36414_o;
  wire [12:0] n36416_o;
  wire [9:0] n36418_o;
  wire [12:0] n36422_o;
  wire [12:0] n36423_o;
  wire n36425_o;
  wire [1:0] n36426_o;
  wire n36428_o;
  wire n36429_o;
  wire [11:0] n36430_o;
  wire [8:0] n36431_o;
  wire [8:0] n36432_o;
  wire [2:0] n36433_o;
  wire [2:0] n36434_o;
  wire [2:0] n36435_o;
  wire n36437_o;
  wire [1:0] n36438_o;
  wire n36440_o;
  wire n36441_o;
  wire n36443_o;
  wire n36444_o;
  wire n36446_o;
  wire [4:0] n36447_o;
  wire [8:0] n36448_o;
  wire [4:0] n36449_o;
  wire [5:0] n36451_o;
  wire [2:0] n36452_o;
  wire [8:0] n36453_o;
  wire [8:0] n36454_o;
  wire [2:0] n36455_o;
  wire [12:0] n36456_o;
  wire n36457_o;
  wire [11:0] n36458_o;
  wire [8:0] n36459_o;
  wire [8:0] n36460_o;
  wire [2:0] n36461_o;
  wire n36463_o;
  wire [4:0] n36464_o;
  wire [8:0] n36465_o;
  wire [4:0] n36466_o;
  wire [5:0] n36468_o;
  wire [2:0] n36469_o;
  wire [8:0] n36470_o;
  wire [8:0] n36471_o;
  wire [2:0] n36472_o;
  wire [11:0] n36473_o;
  wire [11:0] n36474_o;
  wire [11:0] n36475_o;
  wire [11:0] n36476_o;
  wire [11:0] n36477_o;
  wire [11:0] n36480_o;
  wire [11:0] n36481_o;
  wire [1:0] n36497_o;
  wire n36499_o;
  wire n36501_o;
  wire n36502_o;
  wire [2:0] n36503_o;
  wire [12:0] n36515_o;
  wire [12:0] n36516_o;
  wire [12:0] n36517_o;
  wire [9:0] n36519_o;
  wire [12:0] n36523_o;
  wire [12:0] n36524_o;
  wire [12:0] n36526_o;
  wire [9:0] n36528_o;
  wire [12:0] n36532_o;
  wire [12:0] n36533_o;
  wire n36535_o;
  wire [1:0] n36536_o;
  wire n36538_o;
  wire n36539_o;
  wire [11:0] n36540_o;
  wire [8:0] n36541_o;
  wire [8:0] n36542_o;
  wire [2:0] n36543_o;
  wire [2:0] n36544_o;
  wire [2:0] n36545_o;
  wire n36547_o;
  wire [1:0] n36548_o;
  wire n36550_o;
  wire n36551_o;
  wire n36553_o;
  wire n36554_o;
  wire n36556_o;
  wire [4:0] n36557_o;
  wire [8:0] n36558_o;
  wire [4:0] n36559_o;
  wire [5:0] n36561_o;
  wire [2:0] n36562_o;
  wire [8:0] n36563_o;
  wire [8:0] n36564_o;
  wire [2:0] n36565_o;
  wire [12:0] n36566_o;
  wire n36567_o;
  wire [11:0] n36568_o;
  wire [8:0] n36569_o;
  wire [8:0] n36570_o;
  wire [2:0] n36571_o;
  wire n36573_o;
  wire [4:0] n36574_o;
  wire [8:0] n36575_o;
  wire [4:0] n36576_o;
  wire [5:0] n36578_o;
  wire [2:0] n36579_o;
  wire [8:0] n36580_o;
  wire [8:0] n36581_o;
  wire [2:0] n36582_o;
  wire [11:0] n36583_o;
  wire [11:0] n36584_o;
  wire [11:0] n36585_o;
  wire [11:0] n36586_o;
  wire [11:0] n36587_o;
  wire [11:0] n36590_o;
  wire [11:0] n36591_o;
  wire [1:0] n36607_o;
  wire n36609_o;
  wire n36611_o;
  wire n36612_o;
  wire [2:0] n36613_o;
  wire [12:0] n36625_o;
  wire [12:0] n36626_o;
  wire [12:0] n36627_o;
  wire [9:0] n36629_o;
  wire [12:0] n36633_o;
  wire [12:0] n36634_o;
  wire [12:0] n36636_o;
  wire [9:0] n36638_o;
  wire [12:0] n36642_o;
  wire [12:0] n36643_o;
  wire n36645_o;
  wire [1:0] n36646_o;
  wire n36648_o;
  wire n36649_o;
  wire [11:0] n36650_o;
  wire [8:0] n36651_o;
  wire [8:0] n36652_o;
  wire [2:0] n36653_o;
  wire [2:0] n36654_o;
  wire [2:0] n36655_o;
  wire n36657_o;
  wire [1:0] n36658_o;
  wire n36660_o;
  wire n36661_o;
  wire n36663_o;
  wire n36664_o;
  wire n36666_o;
  wire [4:0] n36667_o;
  wire [8:0] n36668_o;
  wire [4:0] n36669_o;
  wire [5:0] n36671_o;
  wire [2:0] n36672_o;
  wire [8:0] n36673_o;
  wire [8:0] n36674_o;
  wire [2:0] n36675_o;
  wire [12:0] n36676_o;
  wire n36677_o;
  wire [11:0] n36678_o;
  wire [8:0] n36679_o;
  wire [8:0] n36680_o;
  wire [2:0] n36681_o;
  wire n36683_o;
  wire [4:0] n36684_o;
  wire [8:0] n36685_o;
  wire [4:0] n36686_o;
  wire [5:0] n36688_o;
  wire [2:0] n36689_o;
  wire [8:0] n36690_o;
  wire [8:0] n36691_o;
  wire [2:0] n36692_o;
  wire [11:0] n36693_o;
  wire [11:0] n36694_o;
  wire [11:0] n36695_o;
  wire [11:0] n36696_o;
  wire [11:0] n36697_o;
  wire [11:0] n36700_o;
  wire [11:0] n36701_o;
  wire [1:0] n36717_o;
  wire n36719_o;
  wire n36721_o;
  wire n36722_o;
  wire [2:0] n36723_o;
  wire [12:0] n36735_o;
  wire [12:0] n36736_o;
  wire [12:0] n36737_o;
  wire [9:0] n36739_o;
  wire [12:0] n36743_o;
  wire [12:0] n36744_o;
  wire [12:0] n36746_o;
  wire [9:0] n36748_o;
  wire [12:0] n36752_o;
  wire [12:0] n36753_o;
  wire n36755_o;
  wire [1:0] n36756_o;
  wire n36758_o;
  wire n36759_o;
  wire [11:0] n36760_o;
  wire [8:0] n36761_o;
  wire [8:0] n36762_o;
  wire [2:0] n36763_o;
  wire [2:0] n36764_o;
  wire [2:0] n36765_o;
  wire n36767_o;
  wire [1:0] n36768_o;
  wire n36770_o;
  wire n36771_o;
  wire n36773_o;
  wire n36774_o;
  wire n36776_o;
  wire [4:0] n36777_o;
  wire [8:0] n36778_o;
  wire [4:0] n36779_o;
  wire [5:0] n36781_o;
  wire [2:0] n36782_o;
  wire [8:0] n36783_o;
  wire [8:0] n36784_o;
  wire [2:0] n36785_o;
  wire [12:0] n36786_o;
  wire n36787_o;
  wire [11:0] n36788_o;
  wire [8:0] n36789_o;
  wire [8:0] n36790_o;
  wire [2:0] n36791_o;
  wire n36793_o;
  wire [4:0] n36794_o;
  wire [8:0] n36795_o;
  wire [4:0] n36796_o;
  wire [5:0] n36798_o;
  wire [2:0] n36799_o;
  wire [8:0] n36800_o;
  wire [8:0] n36801_o;
  wire [2:0] n36802_o;
  wire [11:0] n36803_o;
  wire [11:0] n36804_o;
  wire [11:0] n36805_o;
  wire [11:0] n36806_o;
  wire [11:0] n36807_o;
  wire [11:0] n36810_o;
  wire [11:0] n36811_o;
  wire n36818_o;
  wire [11:0] n36820_o;
  wire [6:0] n36821_o;
  wire [7:0] n36822_o;
  wire [3:0] n36824_o;
  wire [7:0] n36825_o;
  wire [6:0] n36826_o;
  wire [7:0] n36827_o;
  wire [7:0] n36828_o;
  wire n36831_o;
  wire n36833_o;
  wire n36835_o;
  wire n36837_o;
  wire n36839_o;
  wire [4:0] n36841_o;
  wire [7:0] n36846_o;
  wire [7:0] n36848_o;
  wire [7:0] n36850_o;
  wire [7:0] n36852_o;
  reg [3:0] n36923_q;
  reg [3:0] n36924_q;
  reg [3:0] n36925_q;
  reg [3:0] n36926_q;
  reg [3:0] n36927_q;
  reg [3:0] n36928_q;
  reg n36930_q;
  reg n36931_q;
  reg [12:0] n36932_q;
  reg [12:0] n36933_q;
  reg [12:0] n36934_q;
  reg n36935_q;
  reg n36936_q;
  reg n36937_q;
  reg n36938_q;
  reg n36940_q;
  reg n36941_q;
  reg n36942_q;
  reg n36943_q;
  reg n36944_q;
  reg n36945_q;
  reg [11:0] n36946_q;
  reg n36947_q;
  reg n36948_q;
  reg n36949_q;
  reg [4:0] n36950_q;
  wire [11:0] n36951_o;
  reg [11:0] n36952_q;
  wire [11:0] n36953_o;
  reg [11:0] n36954_q;
  wire [11:0] n36955_o;
  reg [11:0] n36956_q;
  reg n36957_q;
  reg n36958_q;
  reg n36959_q;
  reg n36960_q;
  reg n36961_q;
  reg n36962_q;
  reg [4:0] n36964_q;
  reg [3:0] n36965_q;
  reg [3:0] n36966_q;
  reg [3:0] n36967_q;
  reg [12:0] n36968_q;
  reg [4:0] n36969_q;
  reg [3:0] n36970_q;
  reg [3:0] n36971_q;
  reg [3:0] n36972_q;
  reg [3:0] n36973_q;
  reg [3:0] n36974_q;
  reg [12:0] n36975_q;
  reg [12:0] n36976_q;
  reg [2:0] n36977_q;
  reg [2:0] n36978_q;
  reg [2:0] n36979_q;
  reg [2:0] n36980_q;
  reg n36982_q;
  reg n36983_q;
  reg n36984_q;
  reg n36985_q;
  reg [4:0] n36987_q;
  reg [103:0] n36988_q;
  reg [12:0] n36989_q;
  reg [12:0] n36990_q;
  reg [12:0] n36991_q;
  reg [12:0] n36992_q;
  reg [12:0] n36993_q;
  reg [12:0] n36994_q;
  reg [7:0] n36995_q;
  reg [7:0] n36996_q;
  reg [7:0] n36997_q;
  reg [7:0] n36998_q;
  reg [7:0] n36999_q;
  reg [7:0] n37000_q;
  reg [7:0] n37001_q;
  reg [7:0] n37002_q;
  reg [7:0] n37003_q;
  reg [12:0] n37004_q;
  wire [12:0] n37005_o;
  wire [12:0] n37006_o;
  wire [12:0] n37007_o;
  wire [12:0] n37008_o;
  wire [1:0] n37009_o;
  reg [12:0] n37010_o;
  wire [12:0] n37011_o;
  wire [12:0] n37012_o;
  wire [12:0] n37013_o;
  wire [12:0] n37014_o;
  wire [1:0] n37015_o;
  reg [12:0] n37016_o;
  wire [12:0] n37017_o;
  wire [12:0] n37018_o;
  wire [12:0] n37019_o;
  wire [12:0] n37020_o;
  wire [1:0] n37021_o;
  reg [12:0] n37022_o;
  wire [12:0] n37023_o;
  wire [12:0] n37024_o;
  wire [12:0] n37025_o;
  wire [12:0] n37026_o;
  wire [1:0] n37027_o;
  reg [12:0] n37028_o;
  wire [12:0] n37029_o;
  wire [12:0] n37030_o;
  wire [12:0] n37031_o;
  wire [12:0] n37032_o;
  wire [1:0] n37033_o;
  reg [12:0] n37034_o;
  wire [12:0] n37035_o;
  wire [12:0] n37036_o;
  wire [12:0] n37037_o;
  wire [12:0] n37038_o;
  wire [1:0] n37039_o;
  reg [12:0] n37040_o;
  wire [12:0] n37041_o;
  wire [12:0] n37042_o;
  wire [12:0] n37043_o;
  wire [12:0] n37044_o;
  wire [1:0] n37045_o;
  reg [12:0] n37046_o;
  wire [12:0] n37047_o;
  wire [12:0] n37048_o;
  wire [12:0] n37049_o;
  wire [12:0] n37050_o;
  wire [1:0] n37051_o;
  reg [12:0] n37052_o;
  wire [12:0] n37053_o;
  wire [12:0] n37054_o;
  wire [12:0] n37055_o;
  wire [12:0] n37056_o;
  wire [12:0] n37057_o;
  wire [12:0] n37058_o;
  wire [12:0] n37059_o;
  wire [12:0] n37060_o;
  wire [1:0] n37061_o;
  reg [12:0] n37062_o;
  wire [1:0] n37063_o;
  reg [12:0] n37064_o;
  wire n37065_o;
  wire [12:0] n37066_o;
  wire [12:0] n37067_o;
  wire [12:0] n37068_o;
  wire [12:0] n37069_o;
  wire [12:0] n37070_o;
  wire [12:0] n37071_o;
  wire [12:0] n37072_o;
  wire [12:0] n37073_o;
  wire [12:0] n37074_o;
  wire [1:0] n37075_o;
  reg [12:0] n37076_o;
  wire [1:0] n37077_o;
  reg [12:0] n37078_o;
  wire n37079_o;
  wire [12:0] n37080_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n36139_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n35996_o;
  assign i_x2_out = n36033_o;
  assign result_waddr_out = n36034_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n36923_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n36924_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n36925_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n36926_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n36927_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n36928_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n36930_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n36931_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n36932_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n36933_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n36934_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n36935_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n36936_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n36937_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n36938_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n36037_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n36940_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n36941_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n36035_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n36942_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n36057_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n36943_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n36065_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n36944_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n36070_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n36945_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n36946_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n36039_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n36040_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n36041_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n36042_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n36043_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n36044_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n36045_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n36046_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n36047_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n36048_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n36049_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n36050_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n36947_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n36948_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n36949_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n36950_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n36952_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n36954_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n36956_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n36481_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n36591_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n36701_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n36811_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n36957_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n36958_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n36959_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n36960_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n36961_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n36962_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n36192_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n36193_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n36194_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n36195_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n36196_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n36964_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n36965_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n36966_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n36967_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n36968_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n36969_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n36970_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n36971_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n36972_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n36973_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n36974_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n36975_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n36976_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n36977_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n36978_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n36979_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n36980_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n36982_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n36983_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n36984_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n36985_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n36987_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n36988_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n36072_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n36073_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n36989_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n36990_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n36991_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n36992_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n36993_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n36994_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n36082_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n36092_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n36102_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n37028_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n37034_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n37040_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n36137_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n36129_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n37052_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n36995_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n36996_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n36997_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n36998_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n36999_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n37000_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n37001_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n37002_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n37003_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n37004_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n35967_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n35969_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n35972_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n35974_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n35976_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n35978_o = imu_x1_parm_rrr == 4'b1000;
  assign n35979_o = {n35978_o, n35976_o, n35974_o, n35972_o, n35969_o, n35967_o};
  assign n35981_o = imu_const_rrr[3:0];
  assign n35983_o = result_r[3:0];
  assign n35984_o = lane_rrr[3:0];
  assign n35985_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n35979_o)
      6'b100000: n35986_o = n35984_o;
      6'b010000: n35986_o = n35983_o;
      6'b001000: n35986_o = 4'b0001;
      6'b000100: n35986_o = instruction_tid_rrr;
      6'b000010: n35986_o = n35981_o;
      6'b000001: n35986_o = 4'b0000;
      default: n35986_o = n35985_o;
    endcase
  assign n35988_o = imu_const_rrr[12:4];
  assign n35990_o = result_r[12:4];
  assign n35991_o = lane_rrr[12:4];
  assign n35992_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n35979_o)
      6'b100000: n35993_o = n35991_o;
      6'b010000: n35993_o = n35990_o;
      6'b001000: n35993_o = 9'b000000000;
      6'b000100: n35993_o = 9'b000000000;
      6'b000010: n35993_o = n35988_o;
      6'b000001: n35993_o = 9'b000000000;
      default: n35993_o = n35992_o;
    endcase
  assign n35996_o = {n35993_o, n35986_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n36004_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n36006_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n36009_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n36011_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n36013_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n36015_o = imu_x2_parm_rrr == 4'b1000;
  assign n36016_o = {n36015_o, n36013_o, n36011_o, n36009_o, n36006_o, n36004_o};
  assign n36018_o = imu_const_rrr[3:0];
  assign n36020_o = result_r[3:0];
  assign n36021_o = lane_rrr[3:0];
  assign n36022_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n36016_o)
      6'b100000: n36023_o = n36021_o;
      6'b010000: n36023_o = n36020_o;
      6'b001000: n36023_o = 4'b0001;
      6'b000100: n36023_o = instruction_tid_rrr;
      6'b000010: n36023_o = n36018_o;
      6'b000001: n36023_o = 4'b0000;
      default: n36023_o = n36022_o;
    endcase
  assign n36025_o = imu_const_rrr[12:4];
  assign n36027_o = result_r[12:4];
  assign n36028_o = lane_rrr[12:4];
  assign n36029_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n36016_o)
      6'b100000: n36030_o = n36028_o;
      6'b010000: n36030_o = n36027_o;
      6'b001000: n36030_o = 9'b000000000;
      6'b000100: n36030_o = 9'b000000000;
      6'b000010: n36030_o = n36025_o;
      6'b000001: n36030_o = 9'b000000000;
      default: n36030_o = n36029_o;
    endcase
  assign n36033_o = {n36030_o, n36023_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n36034_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n36035_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n36036_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n36037_o = instruction_mu_valid_in ? n36036_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n36039_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n36040_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n36041_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n36042_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n36043_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n36044_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n36045_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n36046_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n36047_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n36048_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n36049_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n36050_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n36053_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n36054_o = n36053_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n36055_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n36056_o = n36055_o & n36054_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n36057_o = n36056_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n36061_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n36062_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n36063_o = n36062_o & n36061_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n36064_o = n36063_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n36065_o = n36064_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n36069_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n36070_o = n36069_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n36072_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n36073_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n36074_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n36078_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n36079_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n36080_o = ~n36079_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n36081_o = n36078_o | n36080_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n36082_o = n36081_o ? n37010_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n36084_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n36088_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n36089_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n36090_o = ~n36089_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n36091_o = n36088_o | n36090_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n36092_o = n36091_o ? n37016_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n36094_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n36098_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n36099_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n36100_o = ~n36099_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n36101_o = n36098_o | n36100_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n36102_o = n36101_o ? n37022_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n36104_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n36108_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n36113_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n36121_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n36125_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n36126_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n36127_o = ~n36126_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n36128_o = n36125_o | n36127_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n36129_o = n36128_o ? n37046_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n36131_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n36135_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n36136_o = ~n36135_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n36137_o = n36136_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n36138_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n36139_o = n36138_o ? mu_lane_rrrrrr : n36140_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n36140_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n36143_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n36145_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n36146_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n36147_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n36148_o = ~n36147_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n36149_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n36150_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n36151_o = n36148_o ? n36149_o : n36150_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n36152_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n36153_o = ~n36152_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n36154_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n36155_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n36156_o = n36153_o ? n36154_o : n36155_o;
  assign n36167_o = {n36145_o, n36151_o, n36156_o, n36146_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n36192_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n36193_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n36194_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n36195_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n36196_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n36200_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n36202_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n36206_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n36211_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n36212_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n36214_o = n36212_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n36215_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n36217_o = n36214_o ? n36215_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n36220_o = n36214_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n36222_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n36225_o = n36222_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n36227_o = n36211_o ? n36225_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n36229_o = n36211_o ? n36217_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n36231_o = n36211_o ? n36220_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n36233_o = got_imu_rr ? n36227_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n36235_o = got_imu_rr ? n36229_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n36237_o = got_imu_rr ? n36231_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n36239_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n36387_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n36389_o = n36387_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n36391_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n36392_o = n36389_o | n36391_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n36393_o = mu_x1_parm1[2:0];
  assign n36405_o = {1'b0, mu_x1_parm1};
  assign n36406_o = {10'b0000000000, n36393_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n36407_o = n36392_o ? n36406_o : n36405_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n36409_o = mu_x1_i1_1[9:0];
  assign n36413_o = {n36409_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n36414_o = mu_x1_vector ? n36413_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n36416_o = mu_x1_i0_1 + n36407_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n36418_o = n36416_o[9:0];
  assign n36422_o = {n36418_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36423_o = mu_x1_vector ? n36422_o : n36416_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n36425_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n36426_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n36428_o = n36426_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n36429_o = n36425_o | n36428_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n36430_o = n36423_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n36431_o = n36430_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n36432_o = ~n36431_o;
  assign n36433_o = n36422_o[2:0];
  assign n36434_o = n36416_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36435_o = mu_x1_vector ? n36433_o : n36434_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n36437_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n36438_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n36440_o = n36438_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n36441_o = n36437_o | n36440_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n36443_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n36444_o = n36441_o | n36443_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n36446_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n36447_o = n36423_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n36448_o = {n36447_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n36449_o = n36423_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n36451_o = {1'b0, n36449_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n36452_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n36453_o = {n36451_o, n36452_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n36454_o = n36446_o ? n36448_o : n36453_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n36455_o = n36423_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n36456_o = n36414_o + n36423_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n36457_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n36458_o = n36456_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n36459_o = n36458_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n36460_o = ~n36459_o;
  assign n36461_o = n36456_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n36463_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n36464_o = n36456_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n36465_o = {n36464_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n36466_o = n36456_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n36468_o = {1'b0, n36466_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n36469_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n36470_o = {n36468_o, n36469_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n36471_o = n36463_o ? n36465_o : n36470_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n36472_o = n36456_o[2:0];
  assign n36473_o = {n36471_o, n36472_o};
  assign n36474_o = {n36460_o, n36461_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n36475_o = n36457_o ? n36474_o : n36473_o;
  assign n36476_o = {n36454_o, n36455_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n36477_o = n36444_o ? n36476_o : n36475_o;
  assign n36480_o = {n36432_o, n36435_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n36481_o = n36429_o ? n36480_o : n36477_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n36497_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n36499_o = n36497_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n36501_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n36502_o = n36499_o | n36501_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n36503_o = mu_x2_parm1[2:0];
  assign n36515_o = {1'b0, mu_x2_parm1};
  assign n36516_o = {10'b0000000000, n36503_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n36517_o = n36502_o ? n36516_o : n36515_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n36519_o = mu_x2_i1_1[9:0];
  assign n36523_o = {n36519_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n36524_o = mu_x2_vector ? n36523_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n36526_o = mu_x2_i0_1 + n36517_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n36528_o = n36526_o[9:0];
  assign n36532_o = {n36528_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36533_o = mu_x2_vector ? n36532_o : n36526_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n36535_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n36536_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n36538_o = n36536_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n36539_o = n36535_o | n36538_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n36540_o = n36533_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n36541_o = n36540_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n36542_o = ~n36541_o;
  assign n36543_o = n36532_o[2:0];
  assign n36544_o = n36526_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36545_o = mu_x2_vector ? n36543_o : n36544_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n36547_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n36548_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n36550_o = n36548_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n36551_o = n36547_o | n36550_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n36553_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n36554_o = n36551_o | n36553_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n36556_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n36557_o = n36533_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n36558_o = {n36557_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n36559_o = n36533_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n36561_o = {1'b0, n36559_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n36562_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n36563_o = {n36561_o, n36562_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n36564_o = n36556_o ? n36558_o : n36563_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n36565_o = n36533_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n36566_o = n36524_o + n36533_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n36567_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n36568_o = n36566_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n36569_o = n36568_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n36570_o = ~n36569_o;
  assign n36571_o = n36566_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n36573_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n36574_o = n36566_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n36575_o = {n36574_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n36576_o = n36566_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n36578_o = {1'b0, n36576_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n36579_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n36580_o = {n36578_o, n36579_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n36581_o = n36573_o ? n36575_o : n36580_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n36582_o = n36566_o[2:0];
  assign n36583_o = {n36581_o, n36582_o};
  assign n36584_o = {n36570_o, n36571_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n36585_o = n36567_o ? n36584_o : n36583_o;
  assign n36586_o = {n36564_o, n36565_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n36587_o = n36554_o ? n36586_o : n36585_o;
  assign n36590_o = {n36542_o, n36545_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n36591_o = n36539_o ? n36590_o : n36587_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n36607_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n36609_o = n36607_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n36611_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n36612_o = n36609_o | n36611_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n36613_o = mu_x3_parm1[2:0];
  assign n36625_o = {1'b0, mu_x3_parm1};
  assign n36626_o = {10'b0000000000, n36613_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n36627_o = n36612_o ? n36626_o : n36625_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n36629_o = mu_x3_i1_1[9:0];
  assign n36633_o = {n36629_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n36634_o = mu_x3_vector ? n36633_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n36636_o = mu_x3_i0_1 + n36627_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n36638_o = n36636_o[9:0];
  assign n36642_o = {n36638_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36643_o = mu_x3_vector ? n36642_o : n36636_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n36645_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n36646_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n36648_o = n36646_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n36649_o = n36645_o | n36648_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n36650_o = n36643_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n36651_o = n36650_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n36652_o = ~n36651_o;
  assign n36653_o = n36642_o[2:0];
  assign n36654_o = n36636_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36655_o = mu_x3_vector ? n36653_o : n36654_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n36657_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n36658_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n36660_o = n36658_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n36661_o = n36657_o | n36660_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n36663_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n36664_o = n36661_o | n36663_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n36666_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n36667_o = n36643_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n36668_o = {n36667_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n36669_o = n36643_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n36671_o = {1'b0, n36669_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n36672_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n36673_o = {n36671_o, n36672_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n36674_o = n36666_o ? n36668_o : n36673_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n36675_o = n36643_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n36676_o = n36634_o + n36643_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n36677_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n36678_o = n36676_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n36679_o = n36678_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n36680_o = ~n36679_o;
  assign n36681_o = n36676_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n36683_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n36684_o = n36676_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n36685_o = {n36684_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n36686_o = n36676_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n36688_o = {1'b0, n36686_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n36689_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n36690_o = {n36688_o, n36689_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n36691_o = n36683_o ? n36685_o : n36690_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n36692_o = n36676_o[2:0];
  assign n36693_o = {n36691_o, n36692_o};
  assign n36694_o = {n36680_o, n36681_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n36695_o = n36677_o ? n36694_o : n36693_o;
  assign n36696_o = {n36674_o, n36675_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n36697_o = n36664_o ? n36696_o : n36695_o;
  assign n36700_o = {n36652_o, n36655_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n36701_o = n36649_o ? n36700_o : n36697_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n36717_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n36719_o = n36717_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n36721_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n36722_o = n36719_o | n36721_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n36723_o = mu_y_parm1[2:0];
  assign n36735_o = {1'b0, mu_y_parm1};
  assign n36736_o = {10'b0000000000, n36723_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n36737_o = n36722_o ? n36736_o : n36735_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n36739_o = mu_y_i1_1[9:0];
  assign n36743_o = {n36739_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n36744_o = mu_y_vector ? n36743_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n36746_o = mu_y_i0_1 + n36737_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n36748_o = n36746_o[9:0];
  assign n36752_o = {n36748_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36753_o = mu_y_vector ? n36752_o : n36746_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n36755_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n36756_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n36758_o = n36756_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n36759_o = n36755_o | n36758_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n36760_o = n36753_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n36761_o = n36760_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n36762_o = ~n36761_o;
  assign n36763_o = n36752_o[2:0];
  assign n36764_o = n36746_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n36765_o = mu_y_vector ? n36763_o : n36764_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n36767_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n36768_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n36770_o = n36768_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n36771_o = n36767_o | n36770_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n36773_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n36774_o = n36771_o | n36773_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n36776_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n36777_o = n36753_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n36778_o = {n36777_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n36779_o = n36753_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n36781_o = {1'b0, n36779_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n36782_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n36783_o = {n36781_o, n36782_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n36784_o = n36776_o ? n36778_o : n36783_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n36785_o = n36753_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n36786_o = n36744_o + n36753_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n36787_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n36788_o = n36786_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n36789_o = n36788_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n36790_o = ~n36789_o;
  assign n36791_o = n36786_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n36793_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n36794_o = n36786_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n36795_o = {n36794_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n36796_o = n36786_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n36798_o = {1'b0, n36796_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n36799_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n36800_o = {n36798_o, n36799_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n36801_o = n36793_o ? n36795_o : n36800_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n36802_o = n36786_o[2:0];
  assign n36803_o = {n36801_o, n36802_o};
  assign n36804_o = {n36790_o, n36791_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n36805_o = n36787_o ? n36804_o : n36803_o;
  assign n36806_o = {n36784_o, n36785_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n36807_o = n36774_o ? n36806_o : n36805_o;
  assign n36810_o = {n36762_o, n36765_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n36811_o = n36759_o ? n36810_o : n36807_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n36818_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n36820_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n36821_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n36822_o = {instruction_vm_in, n36821_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n36824_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n36825_o = {n36824_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n36826_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n36827_o = {instruction_vm_in, n36826_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n36828_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36831_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36833_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36835_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36837_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36839_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36841_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36846_o = instruction_tid_valid_in ? n36828_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36848_o = instruction_tid_valid_in ? n36827_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36850_o = instruction_tid_valid_in ? n36825_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n36852_o = instruction_tid_valid_in ? n36822_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36923_q <= 4'b0000;
    else
      n36923_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36924_q <= 4'b0000;
    else
      n36924_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36925_q <= 4'b0000;
    else
      n36925_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36926_q <= 4'b0000;
    else
      n36926_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36927_q <= 4'b0000;
    else
      n36927_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36928_q <= 4'b0000;
    else
      n36928_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36930_q <= 1'b0;
    else
      n36930_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36931_q <= 1'b0;
    else
      n36931_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36932_q <= 13'b0000000000000;
    else
      n36932_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36933_q <= 13'b0000000000000;
    else
      n36933_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36934_q <= 13'b0000000000000;
    else
      n36934_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36935_q <= 1'b0;
    else
      n36935_q <= n36233_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36936_q <= 1'b0;
    else
      n36936_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36937_q <= 1'b0;
    else
      n36937_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36938_q <= 1'b0;
    else
      n36938_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36940_q <= 1'b0;
    else
      n36940_q <= n36831_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36941_q <= 1'b0;
    else
      n36941_q <= n36833_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36942_q <= 1'b0;
    else
      n36942_q <= n36835_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36943_q <= 1'b0;
    else
      n36943_q <= n36837_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36944_q <= 1'b0;
    else
      n36944_q <= n36839_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36945_q <= 1'b0;
    else
      n36945_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36946_q <= 12'b000000000000;
    else
      n36946_q <= n36820_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36947_q <= 1'b0;
    else
      n36947_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36948_q <= 1'b0;
    else
      n36948_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36949_q <= 1'b0;
    else
      n36949_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36950_q <= 5'b00000;
    else
      n36950_q <= n36841_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n36951_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36952_q <= 12'b000000000000;
    else
      n36952_q <= n36951_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n36953_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36954_q <= 12'b000000000000;
    else
      n36954_q <= n36953_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n36955_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36956_q <= 12'b000000000000;
    else
      n36956_q <= n36955_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36957_q <= 1'b0;
    else
      n36957_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36958_q <= 1'b0;
    else
      n36958_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36959_q <= 1'b0;
    else
      n36959_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36960_q <= 1'b0;
    else
      n36960_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36961_q <= 1'b0;
    else
      n36961_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36962_q <= 1'b0;
    else
      n36962_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36964_q <= 5'b00000;
    else
      n36964_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36965_q <= 4'b0000;
    else
      n36965_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36966_q <= 4'b0000;
    else
      n36966_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36967_q <= 4'b0000;
    else
      n36967_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36968_q <= 13'b0000000000000;
    else
      n36968_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36969_q <= 5'b00000;
    else
      n36969_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36970_q <= 4'b0000;
    else
      n36970_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36971_q <= 4'b0000;
    else
      n36971_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36972_q <= 4'b0000;
    else
      n36972_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36973_q <= 4'b0000;
    else
      n36973_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36974_q <= 4'b0000;
    else
      n36974_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36975_q <= 13'b0000000000000;
    else
      n36975_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36976_q <= 13'b0000000000000;
    else
      n36976_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36977_q <= 3'b000;
    else
      n36977_q <= n36235_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36978_q <= 3'b000;
    else
      n36978_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36979_q <= 3'b000;
    else
      n36979_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36980_q <= 3'b000;
    else
      n36980_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36982_q <= 1'b0;
    else
      n36982_q <= n36237_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36983_q <= 1'b0;
    else
      n36983_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36984_q <= 1'b0;
    else
      n36984_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36985_q <= 1'b0;
    else
      n36985_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36987_q <= 5'b00000;
    else
      n36987_q <= n36239_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n36143_o)
    if (n36143_o)
      n36988_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n36988_q <= n36167_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36989_q <= 13'b0000000000000;
    else
      n36989_q <= n37066_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36990_q <= 13'b0000000000000;
    else
      n36990_q <= n37080_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36991_q <= 13'b0000000000000;
    else
      n36991_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36992_q <= 13'b0000000000000;
    else
      n36992_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36993_q <= 13'b0000000000000;
    else
      n36993_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n36994_q <= 13'b0000000000000;
    else
      n36994_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36995_q <= 8'b00000000;
    else
      n36995_q <= n36846_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36996_q <= 8'b00000000;
    else
      n36996_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36997_q <= 8'b00000000;
    else
      n36997_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36998_q <= 8'b00000000;
    else
      n36998_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n36999_q <= 8'b00000000;
    else
      n36999_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n37000_q <= 8'b00000000;
    else
      n37000_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n37001_q <= 8'b00000000;
    else
      n37001_q <= n36848_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n37002_q <= 8'b00000000;
    else
      n37002_q <= n36850_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n36818_o)
    if (n36818_o)
      n37003_q <= 8'b00000000;
    else
      n37003_q <= n36852_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n36200_o)
    if (n36200_o)
      n37004_q <= 13'b0000000000000;
    else
      n37004_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n37005_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n37006_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n37007_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n37008_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n37009_o = n36074_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n37009_o)
      2'b00: n37010_o = n37005_o;
      2'b01: n37010_o = n37006_o;
      2'b10: n37010_o = n37007_o;
      2'b11: n37010_o = n37008_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n37011_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n37012_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n37013_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n37014_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n37015_o = n36084_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n37015_o)
      2'b00: n37016_o = n37011_o;
      2'b01: n37016_o = n37012_o;
      2'b10: n37016_o = n37013_o;
      2'b11: n37016_o = n37014_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n37017_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n37018_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n37019_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n37020_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n37021_o = n36094_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n37021_o)
      2'b00: n37022_o = n37017_o;
      2'b01: n37022_o = n37018_o;
      2'b10: n37022_o = n37019_o;
      2'b11: n37022_o = n37020_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n37023_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n37024_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n37025_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n37026_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n37027_o = n36104_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n37027_o)
      2'b00: n37028_o = n37023_o;
      2'b01: n37028_o = n37024_o;
      2'b10: n37028_o = n37025_o;
      2'b11: n37028_o = n37026_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n37029_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n37030_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n37031_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n37032_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n37033_o = n36108_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n37033_o)
      2'b00: n37034_o = n37029_o;
      2'b01: n37034_o = n37030_o;
      2'b10: n37034_o = n37031_o;
      2'b11: n37034_o = n37032_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n37035_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n37036_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n37037_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n37038_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n37039_o = n36113_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n37039_o)
      2'b00: n37040_o = n37035_o;
      2'b01: n37040_o = n37036_o;
      2'b10: n37040_o = n37037_o;
      2'b11: n37040_o = n37038_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n37041_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n37042_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n37043_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n37044_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n37045_o = n36121_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n37045_o)
      2'b00: n37046_o = n37041_o;
      2'b01: n37046_o = n37042_o;
      2'b10: n37046_o = n37043_o;
      2'b11: n37046_o = n37044_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n37047_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n37048_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n37049_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n37050_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n37051_o = n36131_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n37051_o)
      2'b00: n37052_o = n37047_o;
      2'b01: n37052_o = n37048_o;
      2'b10: n37052_o = n37049_o;
      2'b11: n37052_o = n37050_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n37053_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n37054_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n37055_o = iregisters_r[38:26];
  assign n37056_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n37057_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n37058_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n37059_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n37060_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n37061_o = n36202_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n37061_o)
      2'b00: n37062_o = n37053_o;
      2'b01: n37062_o = n37054_o;
      2'b10: n37062_o = n37055_o;
      2'b11: n37062_o = n37056_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n37063_o = n36202_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n37063_o)
      2'b00: n37064_o = n37057_o;
      2'b01: n37064_o = n37058_o;
      2'b10: n37064_o = n37059_o;
      2'b11: n37064_o = n37060_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n37065_o = n36202_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n37066_o = n37065_o ? n37064_o : n37062_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n37067_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n37068_o = iregisters_r[25:13];
  assign n37069_o = iregisters_r[38:26];
  assign n37070_o = iregisters_r[51:39];
  assign n37071_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n37072_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n37073_o = iregisters_r[90:78];
  assign n37074_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n37075_o = n36206_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n37075_o)
      2'b00: n37076_o = n37067_o;
      2'b01: n37076_o = n37068_o;
      2'b10: n37076_o = n37069_o;
      2'b11: n37076_o = n37070_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n37077_o = n36206_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n37077_o)
      2'b00: n37078_o = n37071_o;
      2'b01: n37078_o = n37072_o;
      2'b10: n37078_o = n37073_o;
      2'b11: n37078_o = n37074_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n37079_o = n36206_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n37080_o = n37079_o ? n37078_o : n37076_o;
endmodule

module instr_dispatch2
  (input  clock_in,
   input  reset_in,
   input  [4:0] opcode_in,
   input  [3:0] instruction_tid_in,
   input  xreg_in,
   input  flag_in,
   input  wren_in,
   input  en_in,
   input  vm_in,
   input  [11:0] x1_addr1_in,
   input  [11:0] x2_addr1_in,
   input  [11:0] y_addr1_in,
   input  [7:0] result_addr1_in,
   input  x1_vector_in,
   input  x2_vector_in,
   input  y_vector_in,
   input  [7:0] vector_lane_in,
   input  x1_c1_en_in,
   input  [11:0] x1_c1_in,
   input  [95:0] rd_x1_data_in,
   input  [95:0] rd_x2_data_in,
   input  [95:0] mu_y_in,
   output rd_en_out,
   output rd_vm_out,
   output [11:0] rd_x1_addr_out,
   output [11:0] rd_x2_addr_out,
   output rd_x1_vector_out,
   output rd_x2_vector_out,
   output wr_xreg_out,
   output wr_flag_out,
   output wr_xreg_flag_out,
   output wr_en_out,
   output wr_vm_out,
   output wr_vector_out,
   output [11:0] wr_addr_out,
   output [7:0] wr_result_addr_out,
   output [95:0] wr_data_out,
   output [7:0] wr_lane_out,
   output [95:0] mu_x1_out,
   output [95:0] mu_x2_out,
   output [11:0] mu_x_scalar_out,
   output [4:0] mu_opcode_out,
   output [3:0] mu_tid_out);
  wire mu_req;
  wire [4:0] mu_opcode_r;
  wire [4:0] mu_opcode_rr;
  wire [3:0] mu_tid_r;
  wire [3:0] mu_tid_rr;
  wire wr_en_delay;
  wire wr_en_delay_r;
  wire wr_xreg_delay;
  wire wr_xreg_delay_r;
  wire wr_flag_delay;
  wire wr_flag_delay_r;
  wire wr_vm_delay;
  wire wr_vm_delay_r;
  wire [11:0] wr_addr_delay;
  wire [11:0] wr_addr_delay_r;
  wire [7:0] wr_result_addr_delay;
  wire [7:0] wr_result_addr_delay_r;
  wire [7:0] vector_lane_delay;
  wire [7:0] vector_lane_delay_r;
  wire wr_vector_delay;
  wire wr_vector_delay_r;
  wire wr_en;
  wire wr_xreg;
  wire wr_flag;
  wire wr_vm;
  wire x1_c1_en_r;
  wire x1_c1_en_rr;
  wire [11:0] x1_c1_r;
  wire [11:0] x1_c1_rr;
  wire y_vector;
  wire wr_xreg_flag_r;
  wire n35801_o;
  wire n35802_o;
  wire n35803_o;
  wire n35804_o;
  wire n35807_o;
  wire n35808_o;
  wire n35809_o;
  wire n35812_o;
  wire n35813_o;
  wire n35815_o;
  wire n35816_o;
  wire wr_vector_fifo_i_n35817;
  localparam n35818_o = 1'b1;
  wire wr_vector_fifo_i_out_out;
  wire [7:0] wr_vector_lane_fifo_i_n35821;
  localparam n35822_o = 1'b1;
  wire [7:0] wr_vector_lane_fifo_i_out_out;
  wire [11:0] wr_addr_fifo_i_n35825;
  localparam n35826_o = 1'b1;
  wire [11:0] wr_addr_fifo_i_out_out;
  wire [7:0] wr_result_addr_fifo_i_n35829;
  localparam n35830_o = 1'b1;
  wire [7:0] wr_result_addr_fifo_i_out_out;
  wire wr_flag_fifo_i_n35833;
  localparam n35834_o = 1'b1;
  wire wr_flag_fifo_i_out_out;
  wire wr_vm_fifo_i_n35837;
  localparam n35838_o = 1'b1;
  wire wr_vm_fifo_i_out_out;
  wire wr_xreg_fifo_i_n35841;
  localparam n35842_o = 1'b1;
  wire wr_xreg_fifo_i_out_out;
  wire wr_en_fifo_i_n35845;
  localparam n35846_o = 1'b1;
  wire wr_en_fifo_i_out_out;
  wire n35851_o;
  wire n35852_o;
  wire [11:0] n35854_o;
  wire [11:0] n35855_o;
  wire n35858_o;
  wire n35860_o;
  reg [4:0] n35913_q;
  reg [4:0] n35914_q;
  reg [3:0] n35915_q;
  reg [3:0] n35916_q;
  reg n35917_q;
  reg n35918_q;
  reg n35919_q;
  reg n35920_q;
  reg [11:0] n35921_q;
  reg [7:0] n35922_q;
  reg [7:0] n35923_q;
  reg n35924_q;
  reg n35925_q;
  reg n35926_q;
  reg [11:0] n35927_q;
  reg [11:0] n35928_q;
  reg n35929_q;
  assign rd_en_out = en_in;
  assign rd_vm_out = vm_in;
  assign rd_x1_addr_out = x1_addr1_in;
  assign rd_x2_addr_out = x2_addr1_in;
  assign rd_x1_vector_out = x1_vector_in;
  assign rd_x2_vector_out = x2_vector_in;
  assign wr_xreg_out = wr_xreg_delay_r;
  assign wr_flag_out = wr_flag_delay_r;
  assign wr_xreg_flag_out = wr_xreg_flag_r;
  assign wr_en_out = wr_en_delay_r;
  assign wr_vm_out = wr_vm_delay_r;
  assign wr_vector_out = wr_vector_delay_r;
  assign wr_addr_out = wr_addr_delay_r;
  assign wr_result_addr_out = wr_result_addr_delay_r;
  assign wr_data_out = mu_y_in;
  assign wr_lane_out = vector_lane_delay_r;
  assign mu_x1_out = rd_x1_data_in;
  assign mu_x2_out = rd_x2_data_in;
  assign mu_x_scalar_out = n35854_o;
  assign mu_opcode_out = mu_opcode_rr;
  assign mu_tid_out = mu_tid_rr;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:92:8  */
  assign mu_req = n35852_o; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:93:8  */
  assign mu_opcode_r = n35913_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:94:8  */
  assign mu_opcode_rr = n35914_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:95:8  */
  assign mu_tid_r = n35915_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:96:8  */
  assign mu_tid_rr = n35916_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:97:8  */
  assign wr_en_delay = wr_en_fifo_i_n35845; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:98:8  */
  assign wr_en_delay_r = n35917_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:99:8  */
  assign wr_xreg_delay = wr_xreg_fifo_i_n35841; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:100:8  */
  assign wr_xreg_delay_r = n35918_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:101:8  */
  assign wr_flag_delay = wr_flag_fifo_i_n35833; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:102:8  */
  assign wr_flag_delay_r = n35919_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:103:8  */
  assign wr_vm_delay = wr_vm_fifo_i_n35837; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:104:8  */
  assign wr_vm_delay_r = n35920_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:105:8  */
  assign wr_addr_delay = wr_addr_fifo_i_n35825; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:106:8  */
  assign wr_addr_delay_r = n35921_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:107:8  */
  assign wr_result_addr_delay = wr_result_addr_fifo_i_n35829; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:108:8  */
  assign wr_result_addr_delay_r = n35922_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:109:8  */
  assign vector_lane_delay = wr_vector_lane_fifo_i_n35821; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:110:8  */
  assign vector_lane_delay_r = n35923_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:111:8  */
  assign wr_vector_delay = wr_vector_fifo_i_n35817; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:112:8  */
  assign wr_vector_delay_r = n35924_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:113:8  */
  assign wr_en = n35804_o; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:114:8  */
  assign wr_xreg = n35813_o; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:115:8  */
  assign wr_flag = n35809_o; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:116:8  */
  assign wr_vm = vm_in; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:117:8  */
  assign x1_c1_en_r = n35925_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:118:8  */
  assign x1_c1_en_rr = n35926_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:119:8  */
  assign x1_c1_r = n35927_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:120:8  */
  assign x1_c1_rr = n35928_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:121:8  */
  assign y_vector = n35816_o; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:122:8  */
  assign wr_xreg_flag_r = n35929_q; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:126:42  */
  assign n35801_o = ~flag_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:126:31  */
  assign n35802_o = n35801_o & mu_req;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:126:47  */
  assign n35803_o = wren_in & n35802_o;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:126:14  */
  assign n35804_o = n35803_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:128:33  */
  assign n35807_o = flag_in & mu_req;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:128:49  */
  assign n35808_o = wren_in & n35807_o;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:128:16  */
  assign n35809_o = n35808_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:130:33  */
  assign n35812_o = xreg_in & mu_req;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:130:16  */
  assign n35813_o = n35812_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:134:27  */
  assign n35815_o = x1_vector_in | x2_vector_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:134:44  */
  assign n35816_o = wr_flag ? n35815_o : y_vector_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:137:89  */
  assign wr_vector_fifo_i_n35817 = wr_vector_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:136:1  */
  delay_6 wr_vector_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(y_vector),
    .enable_in(n35818_o),
    .out_out(wr_vector_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:140:95  */
  assign wr_vector_lane_fifo_i_n35821 = wr_vector_lane_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:139:1  */
  delayv_8_1 wr_vector_lane_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(vector_lane_in),
    .enable_in(n35822_o),
    .out_out(wr_vector_lane_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:143:91  */
  assign wr_addr_fifo_i_n35825 = wr_addr_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:142:1  */
  delayv_12_6 wr_addr_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(y_addr1_in),
    .enable_in(n35826_o),
    .out_out(wr_addr_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:146:96  */
  assign wr_result_addr_fifo_i_n35829 = wr_result_addr_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:145:1  */
  delayv_8_6 wr_result_addr_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(result_addr1_in),
    .enable_in(n35830_o),
    .out_out(wr_result_addr_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:149:88  */
  assign wr_flag_fifo_i_n35833 = wr_flag_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:148:1  */
  delay_6 wr_flag_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_flag),
    .enable_in(n35834_o),
    .out_out(wr_flag_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:152:86  */
  assign wr_vm_fifo_i_n35837 = wr_vm_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:151:1  */
  delay_6 wr_vm_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_vm),
    .enable_in(n35838_o),
    .out_out(wr_vm_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:155:88  */
  assign wr_xreg_fifo_i_n35841 = wr_xreg_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:154:1  */
  delay_6 wr_xreg_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_xreg),
    .enable_in(n35842_o),
    .out_out(wr_xreg_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:158:86  */
  assign wr_en_fifo_i_n35845 = wr_en_fifo_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_dispatch2.vhd:157:1  */
  delay_6 wr_en_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_en),
    .enable_in(n35846_o),
    .out_out(wr_en_fifo_i_out_out));
  /* ../../HW/src/pcore/instr_dispatch2.vhd:160:30  */
  assign n35851_o = opcode_in == 5'b00000;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:160:15  */
  assign n35852_o = n35851_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:197:29  */
  assign n35854_o = x1_c1_en_rr ? x1_c1_rr : n35855_o;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:197:68  */
  assign n35855_o = rd_x1_data_in[11:0];
  /* ../../HW/src/pcore/instr_dispatch2.vhd:203:16  */
  assign n35858_o = ~reset_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:239:45  */
  assign n35860_o = wr_flag_delay | wr_xreg_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35913_q <= 5'b00000;
    else
      n35913_q <= opcode_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35914_q <= 5'b00000;
    else
      n35914_q <= mu_opcode_r;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35915_q <= 4'b0000;
    else
      n35915_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35916_q <= 4'b0000;
    else
      n35916_q <= mu_tid_r;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35917_q <= 1'b0;
    else
      n35917_q <= wr_en_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35918_q <= 1'b0;
    else
      n35918_q <= wr_xreg_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35919_q <= 1'b0;
    else
      n35919_q <= wr_flag_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35920_q <= 1'b0;
    else
      n35920_q <= wr_vm_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35921_q <= 12'b000000000000;
    else
      n35921_q <= wr_addr_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35922_q <= 8'b00000000;
    else
      n35922_q <= wr_result_addr_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35923_q <= 8'b00000000;
    else
      n35923_q <= vector_lane_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35924_q <= 1'b0;
    else
      n35924_q <= wr_vector_delay;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35925_q <= 1'b0;
    else
      n35925_q <= x1_c1_en_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35926_q <= 1'b0;
    else
      n35926_q <= x1_c1_en_r;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35927_q <= 12'b000000000000;
    else
      n35927_q <= x1_c1_in;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35928_q <= 12'b000000000000;
    else
      n35928_q <= x1_c1_r;
  /* ../../HW/src/pcore/instr_dispatch2.vhd:222:9  */
  always @(posedge clock_in or posedge n35858_o)
    if (n35858_o)
      n35929_q <= 1'b0;
    else
      n35929_q <= n35860_o;
endmodule

module instr_decoder2_0_0
  (input  clock_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  [3:0] instruction_tid_in,
   input  instruction_tid_valid_in,
   input  instruction_vm_in,
   input  [1:0] instruction_data_model_in,
   input  instruction_pre_pre_vm_in,
   input  [1:0] instruction_pre_pre_data_model_in,
   input  [3:0] instruction_pre_tid_in,
   input  instruction_pre_tid_valid_in,
   input  [3:0] instruction_pre_pre_tid_in,
   input  instruction_pre_pre_tid_valid_in,
   input  [27:0] instruction_pre_iregister_auto_in,
   input  [103:0] i_rd_data_in,
   input  [12:0] lane_in,
   input  [12:0] i_y_in,
   input  [12:0] result_in,
   output [4:0] opcode1_out,
   output en1_out,
   output [3:0] instruction_tid_out,
   output xreg1_out,
   output flag1_out,
   output wren_out,
   output vm_out,
   output [11:0] x1_addr1_out,
   output [11:0] x2_addr1_out,
   output [11:0] y_addr1_out,
   output x1_vector_out,
   output x2_vector_out,
   output y_vector_out,
   output [7:0] vector_lane_out,
   output x1_c1_en_out,
   output [11:0] x1_c1_out,
   output i_rd_en_out,
   output i_rd_vm_out,
   output [3:0] i_rd_tid_out,
   output [3:0] i_wr_tid_out,
   output i_wr_en_out,
   output i_wr_vm_out,
   output [2:0] i_wr_addr_out,
   output [12:0] i_wr_data_out,
   output wr_lane_out,
   output [4:0] i_opcode_out,
   output [12:0] i_x1_out,
   output [12:0] i_x2_out,
   output [7:0] result_waddr_out,
   output [7:0] result_raddr_out);
  wire [3:0] instruction_tid_r;
  wire [3:0] instruction_tid_rr;
  wire [3:0] instruction_tid_rrr;
  wire [3:0] instruction_tid_rrrr;
  wire [3:0] instruction_tid_rrrrr;
  wire [3:0] instruction_tid_rrrrrr;
  wire got_imu;
  wire got_imu_r;
  wire got_imu_rr;
  wire [12:0] lane_r;
  wire [12:0] lane_rr;
  wire [12:0] lane_rrr;
  wire imu_lane_valid_r;
  wire imu_lane_valid_rr;
  wire imu_lane_valid_rrr;
  wire imu_lane_valid_rrrr;
  wire [4:0] mu_opcode1;
  wire mu_en1_r;
  wire mu_vm_r;
  wire mu_xreg1;
  wire mu_xreg1_r;
  wire mu_flag1;
  wire mu_flag1_r;
  wire mu_wren;
  wire mu_wren_r;
  wire mu_x1_c1_en;
  wire mu_x1_c1_en_r;
  wire [11:0] mu_x1_c1_r;
  wire [11:0] mu_x1_parm1;
  wire [11:0] mu_x2_parm1;
  wire [11:0] mu_x3_parm1;
  wire [11:0] mu_y_parm1;
  wire [3:0] mu_x1_attr1;
  wire [3:0] mu_x2_attr1;
  wire [3:0] mu_x3_attr1;
  wire [3:0] mu_y_attr1;
  wire mu_x1_vector;
  wire mu_x2_vector;
  wire mu_x3_vector;
  wire mu_y_vector;
  wire mu_x1_vector_r;
  wire mu_x2_vector_r;
  wire mu_y_vector_r;
  wire [4:0] mu_opcode1_r;
  wire [11:0] mu_x1_addr1_r;
  wire [11:0] mu_x2_addr1_r;
  wire [11:0] mu_y_addr1_r;
  wire [11:0] mu_x1_addr1;
  wire [11:0] mu_x2_addr1;
  wire [11:0] mu_x3_addr1;
  wire [11:0] mu_y_addr1;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire vm_rrrrr;
  wire vm_rrrrrr;
  wire [4:0] imu_opcode;
  wire [3:0] imu_x1_parm;
  wire [3:0] imu_x2_parm;
  wire [3:0] imu_y_parm;
  wire [12:0] imu_const;
  wire [4:0] imu_opcode_r;
  wire [3:0] imu_x1_parm_r;
  wire [3:0] imu_x2_parm_r;
  wire [3:0] imu_y_parm_r;
  wire [12:0] imu_const_r;
  wire [4:0] imu_opcode_rr;
  wire [3:0] imu_x1_parm_rr;
  wire [3:0] imu_x2_parm_rr;
  wire [3:0] imu_y_parm_rr;
  wire [3:0] imu_x1_parm_rrr;
  wire [3:0] imu_x2_parm_rrr;
  wire [12:0] imu_const_rr;
  wire [12:0] imu_const_rrr;
  wire [2:0] imu_y_r;
  wire [2:0] imu_y_rr;
  wire [2:0] imu_y_rrr;
  wire [2:0] imu_y_rrrr;
  wire imu_y_valid_r;
  wire imu_y_valid_rr;
  wire imu_y_valid_rrr;
  wire imu_y_valid_rrrr;
  wire [4:0] imu_oc_r;
  wire [103:0] iregisters_r;
  wire [51:0] iregisters_lo;
  wire [51:0] iregisters_hi;
  wire [12:0] imu_x1_ireg_r;
  wire [12:0] imu_x2_ireg_r;
  wire [12:0] imu_x1_ireg_rr;
  wire [12:0] imu_x2_ireg_rr;
  wire [12:0] imu_x1_ireg_rrr;
  wire [12:0] imu_x2_ireg_rrr;
  wire [12:0] mu_x1_i0_1;
  wire [12:0] mu_x2_i0_1;
  wire [12:0] mu_x3_i0_1;
  wire [12:0] mu_x1_i1_1;
  wire [12:0] mu_x2_i1_1;
  wire [12:0] mu_x3_i1_1;
  wire [12:0] mu_x1_i2_1;
  wire [12:0] mu_x1_i2;
  wire [12:0] mu_y_i0_1;
  wire [12:0] mu_y_i1_1;
  wire [7:0] mu_lane_r;
  wire [7:0] mu_lane_rr;
  wire [7:0] mu_lane_rrr;
  wire [7:0] mu_lane_rrrr;
  wire [7:0] mu_lane_rrrrr;
  wire [7:0] mu_lane_rrrrrr;
  wire [7:0] result_raddr_r;
  wire [7:0] result_waddr_r;
  wire [7:0] xreg_waddr_r;
  wire [12:0] result_r;
  wire n34665_o;
  wire n34667_o;
  wire n34670_o;
  wire n34672_o;
  wire n34674_o;
  wire n34676_o;
  wire [5:0] n34677_o;
  wire [3:0] n34679_o;
  wire [3:0] n34681_o;
  wire [3:0] n34682_o;
  wire [3:0] n34683_o;
  reg [3:0] n34684_o;
  wire [8:0] n34686_o;
  wire [8:0] n34688_o;
  wire [8:0] n34689_o;
  wire [8:0] n34690_o;
  reg [8:0] n34691_o;
  wire [12:0] n34694_o;
  wire n34702_o;
  wire n34704_o;
  wire n34707_o;
  wire n34709_o;
  wire n34711_o;
  wire n34713_o;
  wire [5:0] n34714_o;
  wire [3:0] n34716_o;
  wire [3:0] n34718_o;
  wire [3:0] n34719_o;
  wire [3:0] n34720_o;
  reg [3:0] n34721_o;
  wire [8:0] n34723_o;
  wire [8:0] n34725_o;
  wire [8:0] n34726_o;
  wire [8:0] n34727_o;
  reg [8:0] n34728_o;
  wire [12:0] n34731_o;
  wire [7:0] n34732_o;
  wire n34733_o;
  wire [4:0] n34734_o;
  wire [4:0] n34735_o;
  wire [11:0] n34737_o;
  wire [11:0] n34738_o;
  wire [11:0] n34739_o;
  wire [11:0] n34740_o;
  wire [3:0] n34741_o;
  wire [3:0] n34742_o;
  wire [3:0] n34743_o;
  wire [3:0] n34744_o;
  wire n34745_o;
  wire n34746_o;
  wire n34747_o;
  wire n34748_o;
  wire n34751_o;
  wire n34752_o;
  wire n34753_o;
  wire n34754_o;
  wire n34755_o;
  wire n34759_o;
  wire n34760_o;
  wire n34761_o;
  wire n34762_o;
  wire n34763_o;
  wire n34767_o;
  wire n34768_o;
  wire [51:0] n34770_o;
  wire [51:0] n34771_o;
  wire [1:0] n34772_o;
  wire n34776_o;
  wire n34777_o;
  wire n34778_o;
  wire n34779_o;
  wire [12:0] n34780_o;
  wire [1:0] n34782_o;
  wire n34786_o;
  wire n34787_o;
  wire n34788_o;
  wire n34789_o;
  wire [12:0] n34790_o;
  wire [1:0] n34792_o;
  wire n34796_o;
  wire n34797_o;
  wire n34798_o;
  wire n34799_o;
  wire [12:0] n34800_o;
  wire [1:0] n34802_o;
  wire [1:0] n34806_o;
  wire [1:0] n34811_o;
  wire [1:0] n34819_o;
  wire n34823_o;
  wire n34824_o;
  wire n34825_o;
  wire n34826_o;
  wire [12:0] n34827_o;
  wire [1:0] n34829_o;
  wire n34833_o;
  wire n34834_o;
  wire [12:0] n34835_o;
  wire n34836_o;
  wire [7:0] n34837_o;
  wire [7:0] n34838_o;
  wire n34841_o;
  wire [51:0] n34843_o;
  wire [25:0] n34844_o;
  wire n34845_o;
  wire n34846_o;
  wire [12:0] n34847_o;
  wire [12:0] n34848_o;
  wire [12:0] n34849_o;
  wire n34850_o;
  wire n34851_o;
  wire [12:0] n34852_o;
  wire [12:0] n34853_o;
  wire [12:0] n34854_o;
  wire [103:0] n34865_o;
  wire [4:0] n34890_o;
  wire [3:0] n34891_o;
  wire [3:0] n34892_o;
  wire [3:0] n34893_o;
  wire [12:0] n34894_o;
  wire n34898_o;
  wire [2:0] n34900_o;
  wire [2:0] n34904_o;
  wire n34909_o;
  wire n34910_o;
  wire n34912_o;
  wire [2:0] n34913_o;
  wire [2:0] n34915_o;
  wire n34918_o;
  wire n34920_o;
  wire n34923_o;
  wire n34925_o;
  wire [2:0] n34927_o;
  wire n34929_o;
  wire n34931_o;
  wire [2:0] n34933_o;
  wire n34935_o;
  wire [4:0] n34937_o;
  wire [1:0] n35085_o;
  wire n35087_o;
  wire n35089_o;
  wire n35090_o;
  wire [2:0] n35091_o;
  wire [12:0] n35103_o;
  wire [12:0] n35104_o;
  wire [12:0] n35105_o;
  wire [9:0] n35107_o;
  wire [12:0] n35111_o;
  wire [12:0] n35112_o;
  wire [12:0] n35114_o;
  wire [9:0] n35116_o;
  wire [12:0] n35120_o;
  wire [12:0] n35121_o;
  wire n35123_o;
  wire [1:0] n35124_o;
  wire n35126_o;
  wire n35127_o;
  wire [11:0] n35128_o;
  wire [8:0] n35129_o;
  wire [8:0] n35130_o;
  wire [2:0] n35131_o;
  wire [2:0] n35132_o;
  wire [2:0] n35133_o;
  wire n35135_o;
  wire [1:0] n35136_o;
  wire n35138_o;
  wire n35139_o;
  wire n35141_o;
  wire n35142_o;
  wire n35144_o;
  wire [4:0] n35145_o;
  wire [8:0] n35146_o;
  wire [4:0] n35147_o;
  wire [5:0] n35149_o;
  wire [2:0] n35150_o;
  wire [8:0] n35151_o;
  wire [8:0] n35152_o;
  wire [2:0] n35153_o;
  wire [12:0] n35154_o;
  wire n35155_o;
  wire [11:0] n35156_o;
  wire [8:0] n35157_o;
  wire [8:0] n35158_o;
  wire [2:0] n35159_o;
  wire n35161_o;
  wire [4:0] n35162_o;
  wire [8:0] n35163_o;
  wire [4:0] n35164_o;
  wire [5:0] n35166_o;
  wire [2:0] n35167_o;
  wire [8:0] n35168_o;
  wire [8:0] n35169_o;
  wire [2:0] n35170_o;
  wire [11:0] n35171_o;
  wire [11:0] n35172_o;
  wire [11:0] n35173_o;
  wire [11:0] n35174_o;
  wire [11:0] n35175_o;
  wire [11:0] n35178_o;
  wire [11:0] n35179_o;
  wire [1:0] n35195_o;
  wire n35197_o;
  wire n35199_o;
  wire n35200_o;
  wire [2:0] n35201_o;
  wire [12:0] n35213_o;
  wire [12:0] n35214_o;
  wire [12:0] n35215_o;
  wire [9:0] n35217_o;
  wire [12:0] n35221_o;
  wire [12:0] n35222_o;
  wire [12:0] n35224_o;
  wire [9:0] n35226_o;
  wire [12:0] n35230_o;
  wire [12:0] n35231_o;
  wire n35233_o;
  wire [1:0] n35234_o;
  wire n35236_o;
  wire n35237_o;
  wire [11:0] n35238_o;
  wire [8:0] n35239_o;
  wire [8:0] n35240_o;
  wire [2:0] n35241_o;
  wire [2:0] n35242_o;
  wire [2:0] n35243_o;
  wire n35245_o;
  wire [1:0] n35246_o;
  wire n35248_o;
  wire n35249_o;
  wire n35251_o;
  wire n35252_o;
  wire n35254_o;
  wire [4:0] n35255_o;
  wire [8:0] n35256_o;
  wire [4:0] n35257_o;
  wire [5:0] n35259_o;
  wire [2:0] n35260_o;
  wire [8:0] n35261_o;
  wire [8:0] n35262_o;
  wire [2:0] n35263_o;
  wire [12:0] n35264_o;
  wire n35265_o;
  wire [11:0] n35266_o;
  wire [8:0] n35267_o;
  wire [8:0] n35268_o;
  wire [2:0] n35269_o;
  wire n35271_o;
  wire [4:0] n35272_o;
  wire [8:0] n35273_o;
  wire [4:0] n35274_o;
  wire [5:0] n35276_o;
  wire [2:0] n35277_o;
  wire [8:0] n35278_o;
  wire [8:0] n35279_o;
  wire [2:0] n35280_o;
  wire [11:0] n35281_o;
  wire [11:0] n35282_o;
  wire [11:0] n35283_o;
  wire [11:0] n35284_o;
  wire [11:0] n35285_o;
  wire [11:0] n35288_o;
  wire [11:0] n35289_o;
  wire [1:0] n35305_o;
  wire n35307_o;
  wire n35309_o;
  wire n35310_o;
  wire [2:0] n35311_o;
  wire [12:0] n35323_o;
  wire [12:0] n35324_o;
  wire [12:0] n35325_o;
  wire [9:0] n35327_o;
  wire [12:0] n35331_o;
  wire [12:0] n35332_o;
  wire [12:0] n35334_o;
  wire [9:0] n35336_o;
  wire [12:0] n35340_o;
  wire [12:0] n35341_o;
  wire n35343_o;
  wire [1:0] n35344_o;
  wire n35346_o;
  wire n35347_o;
  wire [11:0] n35348_o;
  wire [8:0] n35349_o;
  wire [8:0] n35350_o;
  wire [2:0] n35351_o;
  wire [2:0] n35352_o;
  wire [2:0] n35353_o;
  wire n35355_o;
  wire [1:0] n35356_o;
  wire n35358_o;
  wire n35359_o;
  wire n35361_o;
  wire n35362_o;
  wire n35364_o;
  wire [4:0] n35365_o;
  wire [8:0] n35366_o;
  wire [4:0] n35367_o;
  wire [5:0] n35369_o;
  wire [2:0] n35370_o;
  wire [8:0] n35371_o;
  wire [8:0] n35372_o;
  wire [2:0] n35373_o;
  wire [12:0] n35374_o;
  wire n35375_o;
  wire [11:0] n35376_o;
  wire [8:0] n35377_o;
  wire [8:0] n35378_o;
  wire [2:0] n35379_o;
  wire n35381_o;
  wire [4:0] n35382_o;
  wire [8:0] n35383_o;
  wire [4:0] n35384_o;
  wire [5:0] n35386_o;
  wire [2:0] n35387_o;
  wire [8:0] n35388_o;
  wire [8:0] n35389_o;
  wire [2:0] n35390_o;
  wire [11:0] n35391_o;
  wire [11:0] n35392_o;
  wire [11:0] n35393_o;
  wire [11:0] n35394_o;
  wire [11:0] n35395_o;
  wire [11:0] n35398_o;
  wire [11:0] n35399_o;
  wire [1:0] n35415_o;
  wire n35417_o;
  wire n35419_o;
  wire n35420_o;
  wire [2:0] n35421_o;
  wire [12:0] n35433_o;
  wire [12:0] n35434_o;
  wire [12:0] n35435_o;
  wire [9:0] n35437_o;
  wire [12:0] n35441_o;
  wire [12:0] n35442_o;
  wire [12:0] n35444_o;
  wire [9:0] n35446_o;
  wire [12:0] n35450_o;
  wire [12:0] n35451_o;
  wire n35453_o;
  wire [1:0] n35454_o;
  wire n35456_o;
  wire n35457_o;
  wire [11:0] n35458_o;
  wire [8:0] n35459_o;
  wire [8:0] n35460_o;
  wire [2:0] n35461_o;
  wire [2:0] n35462_o;
  wire [2:0] n35463_o;
  wire n35465_o;
  wire [1:0] n35466_o;
  wire n35468_o;
  wire n35469_o;
  wire n35471_o;
  wire n35472_o;
  wire n35474_o;
  wire [4:0] n35475_o;
  wire [8:0] n35476_o;
  wire [4:0] n35477_o;
  wire [5:0] n35479_o;
  wire [2:0] n35480_o;
  wire [8:0] n35481_o;
  wire [8:0] n35482_o;
  wire [2:0] n35483_o;
  wire [12:0] n35484_o;
  wire n35485_o;
  wire [11:0] n35486_o;
  wire [8:0] n35487_o;
  wire [8:0] n35488_o;
  wire [2:0] n35489_o;
  wire n35491_o;
  wire [4:0] n35492_o;
  wire [8:0] n35493_o;
  wire [4:0] n35494_o;
  wire [5:0] n35496_o;
  wire [2:0] n35497_o;
  wire [8:0] n35498_o;
  wire [8:0] n35499_o;
  wire [2:0] n35500_o;
  wire [11:0] n35501_o;
  wire [11:0] n35502_o;
  wire [11:0] n35503_o;
  wire [11:0] n35504_o;
  wire [11:0] n35505_o;
  wire [11:0] n35508_o;
  wire [11:0] n35509_o;
  wire n35516_o;
  wire [11:0] n35518_o;
  wire [6:0] n35519_o;
  wire [7:0] n35520_o;
  wire [3:0] n35522_o;
  wire [7:0] n35523_o;
  wire [6:0] n35524_o;
  wire [7:0] n35525_o;
  wire [7:0] n35526_o;
  wire n35529_o;
  wire n35531_o;
  wire n35533_o;
  wire n35535_o;
  wire n35537_o;
  wire [4:0] n35539_o;
  wire [7:0] n35544_o;
  wire [7:0] n35546_o;
  wire [7:0] n35548_o;
  wire [7:0] n35550_o;
  reg [3:0] n35621_q;
  reg [3:0] n35622_q;
  reg [3:0] n35623_q;
  reg [3:0] n35624_q;
  reg [3:0] n35625_q;
  reg [3:0] n35626_q;
  reg n35628_q;
  reg n35629_q;
  reg [12:0] n35630_q;
  reg [12:0] n35631_q;
  reg [12:0] n35632_q;
  reg n35633_q;
  reg n35634_q;
  reg n35635_q;
  reg n35636_q;
  reg n35638_q;
  reg n35639_q;
  reg n35640_q;
  reg n35641_q;
  reg n35642_q;
  reg n35643_q;
  reg [11:0] n35644_q;
  reg n35645_q;
  reg n35646_q;
  reg n35647_q;
  reg [4:0] n35648_q;
  wire [11:0] n35649_o;
  reg [11:0] n35650_q;
  wire [11:0] n35651_o;
  reg [11:0] n35652_q;
  wire [11:0] n35653_o;
  reg [11:0] n35654_q;
  reg n35655_q;
  reg n35656_q;
  reg n35657_q;
  reg n35658_q;
  reg n35659_q;
  reg n35660_q;
  reg [4:0] n35662_q;
  reg [3:0] n35663_q;
  reg [3:0] n35664_q;
  reg [3:0] n35665_q;
  reg [12:0] n35666_q;
  reg [4:0] n35667_q;
  reg [3:0] n35668_q;
  reg [3:0] n35669_q;
  reg [3:0] n35670_q;
  reg [3:0] n35671_q;
  reg [3:0] n35672_q;
  reg [12:0] n35673_q;
  reg [12:0] n35674_q;
  reg [2:0] n35675_q;
  reg [2:0] n35676_q;
  reg [2:0] n35677_q;
  reg [2:0] n35678_q;
  reg n35680_q;
  reg n35681_q;
  reg n35682_q;
  reg n35683_q;
  reg [4:0] n35685_q;
  reg [103:0] n35686_q;
  reg [12:0] n35687_q;
  reg [12:0] n35688_q;
  reg [12:0] n35689_q;
  reg [12:0] n35690_q;
  reg [12:0] n35691_q;
  reg [12:0] n35692_q;
  reg [7:0] n35693_q;
  reg [7:0] n35694_q;
  reg [7:0] n35695_q;
  reg [7:0] n35696_q;
  reg [7:0] n35697_q;
  reg [7:0] n35698_q;
  reg [7:0] n35699_q;
  reg [7:0] n35700_q;
  reg [7:0] n35701_q;
  reg [12:0] n35702_q;
  wire [12:0] n35703_o;
  wire [12:0] n35704_o;
  wire [12:0] n35705_o;
  wire [12:0] n35706_o;
  wire [1:0] n35707_o;
  reg [12:0] n35708_o;
  wire [12:0] n35709_o;
  wire [12:0] n35710_o;
  wire [12:0] n35711_o;
  wire [12:0] n35712_o;
  wire [1:0] n35713_o;
  reg [12:0] n35714_o;
  wire [12:0] n35715_o;
  wire [12:0] n35716_o;
  wire [12:0] n35717_o;
  wire [12:0] n35718_o;
  wire [1:0] n35719_o;
  reg [12:0] n35720_o;
  wire [12:0] n35721_o;
  wire [12:0] n35722_o;
  wire [12:0] n35723_o;
  wire [12:0] n35724_o;
  wire [1:0] n35725_o;
  reg [12:0] n35726_o;
  wire [12:0] n35727_o;
  wire [12:0] n35728_o;
  wire [12:0] n35729_o;
  wire [12:0] n35730_o;
  wire [1:0] n35731_o;
  reg [12:0] n35732_o;
  wire [12:0] n35733_o;
  wire [12:0] n35734_o;
  wire [12:0] n35735_o;
  wire [12:0] n35736_o;
  wire [1:0] n35737_o;
  reg [12:0] n35738_o;
  wire [12:0] n35739_o;
  wire [12:0] n35740_o;
  wire [12:0] n35741_o;
  wire [12:0] n35742_o;
  wire [1:0] n35743_o;
  reg [12:0] n35744_o;
  wire [12:0] n35745_o;
  wire [12:0] n35746_o;
  wire [12:0] n35747_o;
  wire [12:0] n35748_o;
  wire [1:0] n35749_o;
  reg [12:0] n35750_o;
  wire [12:0] n35751_o;
  wire [12:0] n35752_o;
  wire [12:0] n35753_o;
  wire [12:0] n35754_o;
  wire [12:0] n35755_o;
  wire [12:0] n35756_o;
  wire [12:0] n35757_o;
  wire [12:0] n35758_o;
  wire [1:0] n35759_o;
  reg [12:0] n35760_o;
  wire [1:0] n35761_o;
  reg [12:0] n35762_o;
  wire n35763_o;
  wire [12:0] n35764_o;
  wire [12:0] n35765_o;
  wire [12:0] n35766_o;
  wire [12:0] n35767_o;
  wire [12:0] n35768_o;
  wire [12:0] n35769_o;
  wire [12:0] n35770_o;
  wire [12:0] n35771_o;
  wire [12:0] n35772_o;
  wire [1:0] n35773_o;
  reg [12:0] n35774_o;
  wire [1:0] n35775_o;
  reg [12:0] n35776_o;
  wire n35777_o;
  wire [12:0] n35778_o;
  assign opcode1_out = mu_opcode1_r;
  assign en1_out = mu_en1_r;
  assign instruction_tid_out = instruction_tid_r;
  assign xreg1_out = mu_xreg1_r;
  assign flag1_out = mu_flag1_r;
  assign wren_out = mu_wren_r;
  assign vm_out = mu_vm_r;
  assign x1_addr1_out = mu_x1_addr1_r;
  assign x2_addr1_out = mu_x2_addr1_r;
  assign y_addr1_out = mu_y_addr1_r;
  assign x1_vector_out = mu_x1_vector_r;
  assign x2_vector_out = mu_x2_vector_r;
  assign y_vector_out = mu_y_vector_r;
  assign vector_lane_out = n34837_o;
  assign x1_c1_en_out = mu_x1_c1_en_r;
  assign x1_c1_out = mu_x1_c1_r;
  assign i_rd_en_out = instruction_pre_pre_tid_valid_in;
  assign i_rd_vm_out = instruction_pre_pre_vm_in;
  assign i_rd_tid_out = instruction_pre_pre_tid_in;
  assign i_wr_tid_out = instruction_tid_rrrrrr;
  assign i_wr_en_out = imu_y_valid_rrrr;
  assign i_wr_vm_out = vm_rrrrrr;
  assign i_wr_addr_out = imu_y_rrrr;
  assign i_wr_data_out = i_y_in;
  assign wr_lane_out = imu_lane_valid_rrrr;
  assign i_opcode_out = imu_oc_r;
  assign i_x1_out = n34694_o;
  assign i_x2_out = n34731_o;
  assign result_waddr_out = n34732_o;
  assign result_raddr_out = result_raddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:125:8  */
  assign instruction_tid_r = n35621_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:126:8  */
  assign instruction_tid_rr = n35622_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:127:8  */
  assign instruction_tid_rrr = n35623_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:128:8  */
  assign instruction_tid_rrrr = n35624_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:129:8  */
  assign instruction_tid_rrrrr = n35625_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:130:8  */
  assign instruction_tid_rrrrrr = n35626_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:132:8  */
  assign got_imu = instruction_imu_valid_in; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:133:8  */
  assign got_imu_r = n35628_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:134:8  */
  assign got_imu_rr = n35629_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:135:8  */
  assign lane_r = n35630_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:136:8  */
  assign lane_rr = n35631_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:137:8  */
  assign lane_rrr = n35632_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:138:8  */
  assign imu_lane_valid_r = n35633_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:139:8  */
  assign imu_lane_valid_rr = n35634_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:140:8  */
  assign imu_lane_valid_rrr = n35635_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:141:8  */
  assign imu_lane_valid_rrrr = n35636_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:148:8  */
  assign mu_opcode1 = n34735_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:149:8  */
  assign mu_en1_r = n35638_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:150:8  */
  assign mu_vm_r = n35639_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:151:8  */
  assign mu_xreg1 = n34733_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:152:8  */
  assign mu_xreg1_r = n35640_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:153:8  */
  assign mu_flag1 = n34755_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:154:8  */
  assign mu_flag1_r = n35641_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:155:8  */
  assign mu_wren = n34763_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:156:8  */
  assign mu_wren_r = n35642_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:157:8  */
  assign mu_x1_c1_en = n34768_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:158:8  */
  assign mu_x1_c1_en_r = n35643_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:159:8  */
  assign mu_x1_c1_r = n35644_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x1_parm1 = n34737_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x2_parm1 = n34738_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_x3_parm1 = n34739_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:4  */
  assign mu_y_parm1 = n34740_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:164:8  */
  assign mu_x1_attr1 = n34741_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:165:8  */
  assign mu_x2_attr1 = n34742_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:166:8  */
  assign mu_x3_attr1 = n34743_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:167:8  */
  assign mu_y_attr1 = n34744_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:168:8  */
  assign mu_x1_vector = n34745_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:169:8  */
  assign mu_x2_vector = n34746_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:170:8  */
  assign mu_x3_vector = n34747_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:171:8  */
  assign mu_y_vector = n34748_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:172:8  */
  assign mu_x1_vector_r = n35645_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:173:8  */
  assign mu_x2_vector_r = n35646_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:174:8  */
  assign mu_y_vector_r = n35647_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:176:8  */
  assign mu_opcode1_r = n35648_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:177:8  */
  assign mu_x1_addr1_r = n35650_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:178:8  */
  assign mu_x2_addr1_r = n35652_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:179:8  */
  assign mu_y_addr1_r = n35654_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:180:8  */
  assign mu_x1_addr1 = n35179_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:181:8  */
  assign mu_x2_addr1 = n35289_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:182:8  */
  assign mu_x3_addr1 = n35399_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:183:8  */
  assign mu_y_addr1 = n35509_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:185:8  */
  assign vm_r = n35655_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:186:8  */
  assign vm_rr = n35656_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:187:8  */
  assign vm_rrr = n35657_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:188:8  */
  assign vm_rrrr = n35658_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:189:8  */
  assign vm_rrrrr = n35659_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:190:8  */
  assign vm_rrrrrr = n35660_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:197:8  */
  assign imu_opcode = n34890_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:198:8  */
  assign imu_x1_parm = n34891_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:199:8  */
  assign imu_x2_parm = n34892_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:200:8  */
  assign imu_y_parm = n34893_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:201:8  */
  assign imu_const = n34894_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:202:8  */
  assign imu_opcode_r = n35662_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:203:8  */
  assign imu_x1_parm_r = n35663_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:204:8  */
  assign imu_x2_parm_r = n35664_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:205:8  */
  assign imu_y_parm_r = n35665_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:206:8  */
  assign imu_const_r = n35666_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:207:8  */
  assign imu_opcode_rr = n35667_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:208:8  */
  assign imu_x1_parm_rr = n35668_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:209:8  */
  assign imu_x2_parm_rr = n35669_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:210:8  */
  assign imu_y_parm_rr = n35670_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:211:8  */
  assign imu_x1_parm_rrr = n35671_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:212:8  */
  assign imu_x2_parm_rrr = n35672_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:213:8  */
  assign imu_const_rr = n35673_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:214:8  */
  assign imu_const_rrr = n35674_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:215:8  */
  assign imu_y_r = n35675_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:216:8  */
  assign imu_y_rr = n35676_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:217:8  */
  assign imu_y_rrr = n35677_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:218:8  */
  assign imu_y_rrrr = n35678_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:220:8  */
  assign imu_y_valid_r = n35680_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:221:8  */
  assign imu_y_valid_rr = n35681_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:222:8  */
  assign imu_y_valid_rrr = n35682_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:223:8  */
  assign imu_y_valid_rrrr = n35683_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:225:8  */
  assign imu_oc_r = n35685_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:232:8  */
  assign iregisters_r = n35686_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:233:8  */
  assign iregisters_lo = n34770_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:234:8  */
  assign iregisters_hi = n34771_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:236:8  */
  assign imu_x1_ireg_r = n35687_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:237:8  */
  assign imu_x2_ireg_r = n35688_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:238:8  */
  assign imu_x1_ireg_rr = n35689_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:239:8  */
  assign imu_x2_ireg_rr = n35690_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:240:8  */
  assign imu_x1_ireg_rrr = n35691_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:241:8  */
  assign imu_x2_ireg_rrr = n35692_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:243:8  */
  assign mu_x1_i0_1 = n34780_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:244:8  */
  assign mu_x2_i0_1 = n34790_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:245:8  */
  assign mu_x3_i0_1 = n34800_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:246:8  */
  assign mu_x1_i1_1 = n35726_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:247:8  */
  assign mu_x2_i1_1 = n35732_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:248:8  */
  assign mu_x3_i1_1 = 13'b0000000000000; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:249:8  */
  assign mu_x1_i2_1 = n35738_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:251:8  */
  assign mu_x1_i2 = n34835_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:253:8  */
  assign mu_y_i0_1 = n34827_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:254:8  */
  assign mu_y_i1_1 = n35750_o; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:257:8  */
  assign mu_lane_r = n35693_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:258:8  */
  assign mu_lane_rr = n35694_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:259:8  */
  assign mu_lane_rrr = n35695_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:260:8  */
  assign mu_lane_rrrr = n35696_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:261:8  */
  assign mu_lane_rrrrr = n35697_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:262:8  */
  assign mu_lane_rrrrrr = n35698_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:265:8  */
  assign result_raddr_r = n35699_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:266:8  */
  assign result_waddr_r = n35700_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:267:8  */
  assign xreg_waddr_r = n35701_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:269:8  */
  assign result_r = n35702_q; // (signal)
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n34665_o = imu_x1_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n34667_o = imu_x1_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n34670_o = imu_x1_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n34672_o = imu_x1_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n34674_o = imu_x1_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n34676_o = imu_x1_parm_rrr == 4'b1000;
  assign n34677_o = {n34676_o, n34674_o, n34672_o, n34670_o, n34667_o, n34665_o};
  assign n34679_o = imu_const_rrr[3:0];
  assign n34681_o = result_r[3:0];
  assign n34682_o = lane_rrr[3:0];
  assign n34683_o = imu_x1_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n34677_o)
      6'b100000: n34684_o = n34682_o;
      6'b010000: n34684_o = n34681_o;
      6'b001000: n34684_o = 4'b0000;
      6'b000100: n34684_o = instruction_tid_rrr;
      6'b000010: n34684_o = n34679_o;
      6'b000001: n34684_o = 4'b0000;
      default: n34684_o = n34683_o;
    endcase
  assign n34686_o = imu_const_rrr[12:4];
  assign n34688_o = result_r[12:4];
  assign n34689_o = lane_rrr[12:4];
  assign n34690_o = imu_x1_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n34677_o)
      6'b100000: n34691_o = n34689_o;
      6'b010000: n34691_o = n34688_o;
      6'b001000: n34691_o = 9'b000000000;
      6'b000100: n34691_o = 9'b000000000;
      6'b000010: n34691_o = n34686_o;
      6'b000001: n34691_o = 9'b000000000;
      default: n34691_o = n34690_o;
    endcase
  assign n34694_o = {n34691_o, n34684_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:380:5  */
  assign n34702_o = imu_x2_parm_rrr == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:382:5  */
  assign n34704_o = imu_x2_parm_rrr == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:384:5  */
  assign n34707_o = imu_x2_parm_rrr == 4'b1100;
  /* ../../HW/src/pcore/instr_decoder2.vhd:387:5  */
  assign n34709_o = imu_x2_parm_rrr == 4'b1101;
  /* ../../HW/src/pcore/instr_decoder2.vhd:389:5  */
  assign n34711_o = imu_x2_parm_rrr == 4'b1110;
  /* ../../HW/src/pcore/instr_decoder2.vhd:391:5  */
  assign n34713_o = imu_x2_parm_rrr == 4'b1000;
  assign n34714_o = {n34713_o, n34711_o, n34709_o, n34707_o, n34704_o, n34702_o};
  assign n34716_o = imu_const_rrr[3:0];
  assign n34718_o = result_r[3:0];
  assign n34719_o = lane_rrr[3:0];
  assign n34720_o = imu_x2_ireg_rrr[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n34714_o)
      6'b100000: n34721_o = n34719_o;
      6'b010000: n34721_o = n34718_o;
      6'b001000: n34721_o = 4'b0000;
      6'b000100: n34721_o = instruction_tid_rrr;
      6'b000010: n34721_o = n34716_o;
      6'b000001: n34721_o = 4'b0000;
      default: n34721_o = n34720_o;
    endcase
  assign n34723_o = imu_const_rrr[12:4];
  assign n34725_o = result_r[12:4];
  assign n34726_o = lane_rrr[12:4];
  assign n34727_o = imu_x2_ireg_rrr[12:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:379:1  */
  always @*
    case (n34714_o)
      6'b100000: n34728_o = n34726_o;
      6'b010000: n34728_o = n34725_o;
      6'b001000: n34728_o = 9'b000000000;
      6'b000100: n34728_o = 9'b000000000;
      6'b000010: n34728_o = n34723_o;
      6'b000001: n34728_o = 9'b000000000;
      default: n34728_o = n34727_o;
    endcase
  assign n34731_o = {n34728_o, n34721_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:416:34  */
  assign n34732_o = mu_xreg1_r ? xreg_waddr_r : result_waddr_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:419:30  */
  assign n34733_o = instruction_mu_in[74];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:32  */
  assign n34734_o = instruction_mu_in[79:75];
  /* ../../HW/src/pcore/instr_decoder2.vhd:425:87  */
  assign n34735_o = instruction_mu_valid_in ? n34734_o : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:426:33  */
  assign n34737_o = instruction_mu_in[49:38];
  /* ../../HW/src/pcore/instr_decoder2.vhd:427:33  */
  assign n34738_o = instruction_mu_in[32:21];
  /* ../../HW/src/pcore/instr_decoder2.vhd:428:33  */
  assign n34739_o = instruction_mu_in[66:55];
  /* ../../HW/src/pcore/instr_decoder2.vhd:429:32  */
  assign n34740_o = instruction_mu_in[15:4];
  /* ../../HW/src/pcore/instr_decoder2.vhd:430:33  */
  assign n34741_o = instruction_mu_in[37:34];
  /* ../../HW/src/pcore/instr_decoder2.vhd:431:33  */
  assign n34742_o = instruction_mu_in[20:17];
  /* ../../HW/src/pcore/instr_decoder2.vhd:432:33  */
  assign n34743_o = instruction_mu_in[54:51];
  /* ../../HW/src/pcore/instr_decoder2.vhd:433:32  */
  assign n34744_o = instruction_mu_in[3:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:434:34  */
  assign n34745_o = instruction_mu_in[50];
  /* ../../HW/src/pcore/instr_decoder2.vhd:435:34  */
  assign n34746_o = instruction_mu_in[33];
  /* ../../HW/src/pcore/instr_decoder2.vhd:436:34  */
  assign n34747_o = instruction_mu_in[67];
  /* ../../HW/src/pcore/instr_decoder2.vhd:437:33  */
  assign n34748_o = instruction_mu_in[16];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:65  */
  assign n34751_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:51  */
  assign n34752_o = n34751_o & instruction_mu_valid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:87  */
  assign n34753_o = mu_y_parm1[6];
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:73  */
  assign n34754_o = n34753_o & n34752_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:438:17  */
  assign n34755_o = n34754_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:32  */
  assign n34759_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:54  */
  assign n34760_o = mu_y_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:40  */
  assign n34761_o = n34760_o & n34759_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:88  */
  assign n34762_o = n34761_o | mu_xreg1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:439:16  */
  assign n34763_o = n34762_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:37  */
  assign n34767_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:443:20  */
  assign n34768_o = n34767_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:450:30  */
  assign n34770_o = iregisters_r[51:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:453:30  */
  assign n34771_o = iregisters_r[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:60  */
  assign n34772_o = mu_x1_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:92  */
  assign n34776_o = mu_x1_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:114  */
  assign n34777_o = mu_x1_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:117  */
  assign n34778_o = ~n34777_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:100  */
  assign n34779_o = n34776_o | n34778_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:76  */
  assign n34780_o = n34779_o ? n35708_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:60  */
  assign n34782_o = mu_x2_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:92  */
  assign n34786_o = mu_x2_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:114  */
  assign n34787_o = mu_x2_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:117  */
  assign n34788_o = ~n34787_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:100  */
  assign n34789_o = n34786_o | n34788_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:76  */
  assign n34790_o = n34789_o ? n35714_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:60  */
  assign n34792_o = mu_x3_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:92  */
  assign n34796_o = mu_x3_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:114  */
  assign n34797_o = mu_x3_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:117  */
  assign n34798_o = ~n34797_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:100  */
  assign n34799_o = n34796_o | n34798_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:76  */
  assign n34800_o = n34799_o ? n35720_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:60  */
  assign n34802_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:60  */
  assign n34806_o = mu_x2_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:60  */
  assign n34811_o = mu_x1_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:58  */
  assign n34819_o = mu_y_attr1[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:89  */
  assign n34823_o = mu_y_attr1[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:110  */
  assign n34824_o = mu_y_attr1[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:113  */
  assign n34825_o = ~n34824_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:97  */
  assign n34826_o = n34823_o | n34825_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:74  */
  assign n34827_o = n34826_o ? n35744_o : 13'b0000000000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:58  */
  assign n34829_o = mu_y_parm1[4:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:40  */
  assign n34833_o = mu_x1_parm1[5];
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:43  */
  assign n34834_o = ~n34833_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:469:24  */
  assign n34835_o = n34834_o ? mu_x1_i2_1 : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:59  */
  assign n34836_o = ~imu_lane_valid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:35  */
  assign n34837_o = n34836_o ? mu_lane_rrrrrr : n34838_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:481:92  */
  assign n34838_o = i_y_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:497:12  */
  assign n34841_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:520:81  */
  assign n34843_o = i_rd_data_in[103:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:521:88  */
  assign n34844_o = i_rd_data_in[25:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n34845_o = instruction_pre_iregister_auto_in[26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n34846_o = ~n34845_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n34847_o = i_rd_data_in[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n34848_o = instruction_pre_iregister_auto_in[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n34849_o = n34846_o ? n34847_o : n34848_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:48  */
  assign n34850_o = instruction_pre_iregister_auto_in[27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:96  */
  assign n34851_o = ~n34850_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:524:66  */
  assign n34852_o = i_rd_data_in[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:526:87  */
  assign n34853_o = instruction_pre_iregister_auto_in[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:523:12  */
  assign n34854_o = n34851_o ? n34852_o : n34853_o;
  assign n34865_o = {n34843_o, n34849_o, n34854_o, n34844_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:544:33  */
  assign n34890_o = instruction_imu_in[31:27];
  /* ../../HW/src/pcore/instr_decoder2.vhd:545:34  */
  assign n34891_o = instruction_imu_in[26:23];
  /* ../../HW/src/pcore/instr_decoder2.vhd:546:34  */
  assign n34892_o = instruction_imu_in[22:19];
  /* ../../HW/src/pcore/instr_decoder2.vhd:547:33  */
  assign n34893_o = instruction_imu_in[18:15];
  /* ../../HW/src/pcore/instr_decoder2.vhd:548:41  */
  assign n34894_o = instruction_imu_in[14:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:559:12  */
  assign n34898_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:70  */
  assign n34900_o = imu_x1_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:70  */
  assign n34904_o = imu_x2_parm[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:30  */
  assign n34909_o = imu_opcode_rr != 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:42  */
  assign n34910_o = imu_y_parm_rr[3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:98  */
  assign n34912_o = n34910_o == 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:653:54  */
  assign n34913_o = imu_y_parm_rr[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n34915_o = n34912_o ? n34913_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:652:17  */
  assign n34918_o = n34912_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:33  */
  assign n34920_o = imu_y_parm_rr == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:659:17  */
  assign n34923_o = n34920_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n34925_o = n34909_o ? n34923_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n34927_o = n34909_o ? n34915_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:651:13  */
  assign n34929_o = n34909_o ? n34918_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n34931_o = got_imu_rr ? n34925_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n34933_o = got_imu_rr ? n34927_o : 3'b000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n34935_o = got_imu_rr ? n34929_o : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:648:9  */
  assign n34937_o = got_imu_rr ? imu_opcode_rr : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n35085_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n35087_o = n35085_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n35089_o = mu_x1_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n35090_o = n35087_o | n35089_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n35091_o = mu_x1_parm1[2:0];
  assign n35103_o = {1'b0, mu_x1_parm1};
  assign n35104_o = {10'b0000000000, n35091_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n35105_o = n35090_o ? n35104_o : n35103_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n35107_o = mu_x1_i1_1[9:0];
  assign n35111_o = {n35107_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n35112_o = mu_x1_vector ? n35111_o : mu_x1_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n35114_o = mu_x1_i0_1 + n35105_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n35116_o = n35114_o[9:0];
  assign n35120_o = {n35116_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35121_o = mu_x1_vector ? n35120_o : n35114_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n35123_o = mu_x1_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n35124_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n35126_o = n35124_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n35127_o = n35123_o | n35126_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n35128_o = n35121_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n35129_o = n35128_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n35130_o = ~n35129_o;
  assign n35131_o = n35120_o[2:0];
  assign n35132_o = n35114_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35133_o = mu_x1_vector ? n35131_o : n35132_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n35135_o = mu_x1_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n35136_o = mu_x1_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n35138_o = n35136_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n35139_o = n35135_o | n35138_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n35141_o = mu_x1_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n35142_o = n35139_o | n35141_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n35144_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n35145_o = n35121_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n35146_o = {n35145_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n35147_o = n35121_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n35149_o = {1'b0, n35147_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n35150_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n35151_o = {n35149_o, n35150_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n35152_o = n35144_o ? n35146_o : n35151_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n35153_o = n35121_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n35154_o = n35112_o + n35121_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n35155_o = mu_x1_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n35156_o = n35154_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n35157_o = n35156_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n35158_o = ~n35157_o;
  assign n35159_o = n35154_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n35161_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n35162_o = n35154_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n35163_o = {n35162_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n35164_o = n35154_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n35166_o = {1'b0, n35164_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n35167_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n35168_o = {n35166_o, n35167_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n35169_o = n35161_o ? n35163_o : n35168_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n35170_o = n35154_o[2:0];
  assign n35171_o = {n35169_o, n35170_o};
  assign n35172_o = {n35158_o, n35159_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n35173_o = n35155_o ? n35172_o : n35171_o;
  assign n35174_o = {n35152_o, n35153_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n35175_o = n35142_o ? n35174_o : n35173_o;
  assign n35178_o = {n35130_o, n35133_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n35179_o = n35127_o ? n35178_o : n35175_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n35195_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n35197_o = n35195_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n35199_o = mu_x2_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n35200_o = n35197_o | n35199_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n35201_o = mu_x2_parm1[2:0];
  assign n35213_o = {1'b0, mu_x2_parm1};
  assign n35214_o = {10'b0000000000, n35201_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n35215_o = n35200_o ? n35214_o : n35213_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n35217_o = mu_x2_i1_1[9:0];
  assign n35221_o = {n35217_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n35222_o = mu_x2_vector ? n35221_o : mu_x2_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n35224_o = mu_x2_i0_1 + n35215_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n35226_o = n35224_o[9:0];
  assign n35230_o = {n35226_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35231_o = mu_x2_vector ? n35230_o : n35224_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n35233_o = mu_x2_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n35234_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n35236_o = n35234_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n35237_o = n35233_o | n35236_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n35238_o = n35231_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n35239_o = n35238_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n35240_o = ~n35239_o;
  assign n35241_o = n35230_o[2:0];
  assign n35242_o = n35224_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35243_o = mu_x2_vector ? n35241_o : n35242_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n35245_o = mu_x2_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n35246_o = mu_x2_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n35248_o = n35246_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n35249_o = n35245_o | n35248_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n35251_o = mu_x2_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n35252_o = n35249_o | n35251_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n35254_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n35255_o = n35231_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n35256_o = {n35255_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n35257_o = n35231_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n35259_o = {1'b0, n35257_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n35260_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n35261_o = {n35259_o, n35260_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n35262_o = n35254_o ? n35256_o : n35261_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n35263_o = n35231_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n35264_o = n35222_o + n35231_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n35265_o = mu_x2_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n35266_o = n35264_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n35267_o = n35266_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n35268_o = ~n35267_o;
  assign n35269_o = n35264_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n35271_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n35272_o = n35264_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n35273_o = {n35272_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n35274_o = n35264_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n35276_o = {1'b0, n35274_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n35277_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n35278_o = {n35276_o, n35277_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n35279_o = n35271_o ? n35273_o : n35278_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n35280_o = n35264_o[2:0];
  assign n35281_o = {n35279_o, n35280_o};
  assign n35282_o = {n35268_o, n35269_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n35283_o = n35265_o ? n35282_o : n35281_o;
  assign n35284_o = {n35262_o, n35263_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n35285_o = n35252_o ? n35284_o : n35283_o;
  assign n35288_o = {n35240_o, n35243_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n35289_o = n35237_o ? n35288_o : n35285_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n35305_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n35307_o = n35305_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n35309_o = mu_x3_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n35310_o = n35307_o | n35309_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n35311_o = mu_x3_parm1[2:0];
  assign n35323_o = {1'b0, mu_x3_parm1};
  assign n35324_o = {10'b0000000000, n35311_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n35325_o = n35310_o ? n35324_o : n35323_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n35327_o = mu_x3_i1_1[9:0];
  assign n35331_o = {n35327_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n35332_o = mu_x3_vector ? n35331_o : mu_x3_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n35334_o = mu_x3_i0_1 + n35325_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n35336_o = n35334_o[9:0];
  assign n35340_o = {n35336_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35341_o = mu_x3_vector ? n35340_o : n35334_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n35343_o = mu_x3_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n35344_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n35346_o = n35344_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n35347_o = n35343_o | n35346_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n35348_o = n35341_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n35349_o = n35348_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n35350_o = ~n35349_o;
  assign n35351_o = n35340_o[2:0];
  assign n35352_o = n35334_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35353_o = mu_x3_vector ? n35351_o : n35352_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n35355_o = mu_x3_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n35356_o = mu_x3_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n35358_o = n35356_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n35359_o = n35355_o | n35358_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n35361_o = mu_x3_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n35362_o = n35359_o | n35361_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n35364_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n35365_o = n35341_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n35366_o = {n35365_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n35367_o = n35341_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n35369_o = {1'b0, n35367_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n35370_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n35371_o = {n35369_o, n35370_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n35372_o = n35364_o ? n35366_o : n35371_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n35373_o = n35341_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n35374_o = n35332_o + n35341_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n35375_o = mu_x3_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n35376_o = n35374_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n35377_o = n35376_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n35378_o = ~n35377_o;
  assign n35379_o = n35374_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n35381_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n35382_o = n35374_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n35383_o = {n35382_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n35384_o = n35374_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n35386_o = {1'b0, n35384_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n35387_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n35388_o = {n35386_o, n35387_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n35389_o = n35381_o ? n35383_o : n35388_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n35390_o = n35374_o[2:0];
  assign n35391_o = {n35389_o, n35390_o};
  assign n35392_o = {n35378_o, n35379_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n35393_o = n35375_o ? n35392_o : n35391_o;
  assign n35394_o = {n35372_o, n35373_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n35395_o = n35362_o ? n35394_o : n35393_o;
  assign n35398_o = {n35350_o, n35353_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n35399_o = n35347_o ? n35398_o : n35395_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:11  */
  assign n35415_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:23  */
  assign n35417_o = n35415_o == 2'b11;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:39  */
  assign n35419_o = mu_y_attr1 == 4'b1011;
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:29  */
  assign n35420_o = n35417_o | n35419_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:304:44  */
  assign n35421_o = mu_y_parm1[2:0];
  assign n35433_o = {1'b0, mu_y_parm1};
  assign n35434_o = {10'b0000000000, n35421_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:302:1  */
  assign n35435_o = n35420_o ? n35434_o : n35433_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:317:42  */
  assign n35437_o = mu_y_i1_1[9:0];
  assign n35441_o = {n35437_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:316:1  */
  assign n35442_o = mu_y_vector ? n35441_o : mu_y_i1_1;
  /* ../../HW/src/pcore/instr_decoder2.vhd:325:15  */
  assign n35444_o = mu_y_i0_1 + n35435_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:327:43  */
  assign n35446_o = n35444_o[9:0];
  assign n35450_o = {n35446_o, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35451_o = mu_y_vector ? n35450_o : n35444_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:11  */
  assign n35453_o = mu_y_attr1 == 4'b1000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:29  */
  assign n35454_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:41  */
  assign n35456_o = n35454_o == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:19  */
  assign n35457_o = n35453_o | n35456_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:335:70  */
  assign n35458_o = n35451_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:72  */
  assign n35459_o = n35458_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:336:62  */
  assign n35460_o = ~n35459_o;
  assign n35461_o = n35450_o[2:0];
  assign n35462_o = n35444_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:326:1  */
  assign n35463_o = mu_y_vector ? n35461_o : n35462_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:14  */
  assign n35465_o = mu_y_attr1 == 4'b1001;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:32  */
  assign n35466_o = mu_y_attr1[3:2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:44  */
  assign n35468_o = n35466_o == 2'b01;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:22  */
  assign n35469_o = n35465_o | n35468_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:60  */
  assign n35471_o = mu_y_attr1 == 4'b1010;
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:50  */
  assign n35472_o = n35469_o | n35471_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:20  */
  assign n35474_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:86  */
  assign n35475_o = n35451_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:340:130  */
  assign n35476_o = {n35475_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:92  */
  assign n35477_o = n35451_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:68  */
  assign n35479_o = {1'b0, n35477_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:161  */
  assign n35480_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:342:136  */
  assign n35481_o = {n35479_o, n35480_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:339:4  */
  assign n35482_o = n35474_o ? n35476_o : n35481_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:344:63  */
  assign n35483_o = n35451_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:347:23  */
  assign n35484_o = n35442_o + n35451_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:12  */
  assign n35485_o = mu_y_i1_1[12];
  /* ../../HW/src/pcore/instr_decoder2.vhd:350:79  */
  assign n35486_o = n35484_o[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:75  */
  assign n35487_o = n35486_o[11:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:351:65  */
  assign n35488_o = ~n35487_o;
  assign n35489_o = n35484_o[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:23  */
  assign n35491_o = instruction_data_model_in == 2'b00;
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:95  */
  assign n35492_o = n35484_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:354:139  */
  assign n35493_o = {n35492_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:101  */
  assign n35494_o = n35484_o[7:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:71  */
  assign n35496_o = {1'b0, n35494_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:170  */
  assign n35497_o = instruction_tid_in[2:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:356:145  */
  assign n35498_o = {n35496_o, n35497_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:353:7  */
  assign n35499_o = n35491_o ? n35493_o : n35498_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:358:72  */
  assign n35500_o = n35484_o[2:0];
  assign n35501_o = {n35499_o, n35500_o};
  assign n35502_o = {n35488_o, n35489_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:348:4  */
  assign n35503_o = n35485_o ? n35502_o : n35501_o;
  assign n35504_o = {n35482_o, n35483_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:337:1  */
  assign n35505_o = n35472_o ? n35504_o : n35503_o;
  assign n35508_o = {n35460_o, n35463_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:333:1  */
  assign n35509_o = n35457_o ? n35508_o : n35505_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:713:17  */
  assign n35516_o = ~reset_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:744:52  */
  assign n35518_o = mu_x1_i2[11:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:63  */
  assign n35519_o = mu_y_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:748:51  */
  assign n35520_o = {instruction_vm_in, n35519_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:53  */
  assign n35522_o = {instruction_vm_in, 3'b000};
  /* ../../HW/src/pcore/instr_decoder2.vhd:749:114  */
  assign n35523_o = {n35522_o, instruction_tid_in};
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:66  */
  assign n35524_o = mu_x3_addr1[9:3];
  /* ../../HW/src/pcore/instr_decoder2.vhd:754:53  */
  assign n35525_o = {instruction_vm_in, n35524_o};
  /* ../../HW/src/pcore/instr_decoder2.vhd:755:54  */
  assign n35526_o = lane_in[7:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35529_o = instruction_tid_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35531_o = instruction_tid_valid_in ? instruction_vm_in : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35533_o = instruction_tid_valid_in ? mu_xreg1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35535_o = instruction_tid_valid_in ? mu_flag1 : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35537_o = instruction_tid_valid_in ? mu_wren : 1'b0;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35539_o = instruction_tid_valid_in ? mu_opcode1 : 5'b00000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35544_o = instruction_tid_valid_in ? n35526_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35546_o = instruction_tid_valid_in ? n35525_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35548_o = instruction_tid_valid_in ? n35523_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:746:13  */
  assign n35550_o = instruction_tid_valid_in ? n35520_o : 8'b00000000;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35621_q <= 4'b0000;
    else
      n35621_q <= instruction_tid_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35622_q <= 4'b0000;
    else
      n35622_q <= instruction_tid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35623_q <= 4'b0000;
    else
      n35623_q <= instruction_tid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35624_q <= 4'b0000;
    else
      n35624_q <= instruction_tid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35625_q <= 4'b0000;
    else
      n35625_q <= instruction_tid_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35626_q <= 4'b0000;
    else
      n35626_q <= instruction_tid_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35628_q <= 1'b0;
    else
      n35628_q <= got_imu;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35629_q <= 1'b0;
    else
      n35629_q <= got_imu_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35630_q <= 13'b0000000000000;
    else
      n35630_q <= lane_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35631_q <= 13'b0000000000000;
    else
      n35631_q <= lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35632_q <= 13'b0000000000000;
    else
      n35632_q <= lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35633_q <= 1'b0;
    else
      n35633_q <= n34931_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35634_q <= 1'b0;
    else
      n35634_q <= imu_lane_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35635_q <= 1'b0;
    else
      n35635_q <= imu_lane_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35636_q <= 1'b0;
    else
      n35636_q <= imu_lane_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35638_q <= 1'b0;
    else
      n35638_q <= n35529_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35639_q <= 1'b0;
    else
      n35639_q <= n35531_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35640_q <= 1'b0;
    else
      n35640_q <= n35533_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35641_q <= 1'b0;
    else
      n35641_q <= n35535_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35642_q <= 1'b0;
    else
      n35642_q <= n35537_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35643_q <= 1'b0;
    else
      n35643_q <= mu_x1_c1_en;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35644_q <= 12'b000000000000;
    else
      n35644_q <= n35518_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35645_q <= 1'b0;
    else
      n35645_q <= mu_x1_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35646_q <= 1'b0;
    else
      n35646_q <= mu_x2_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35647_q <= 1'b0;
    else
      n35647_q <= mu_y_vector;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35648_q <= 5'b00000;
    else
      n35648_q <= n35539_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n35649_o = instruction_tid_valid_in ? mu_x1_addr1 : mu_x1_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35650_q <= 12'b000000000000;
    else
      n35650_q <= n35649_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n35651_o = instruction_tid_valid_in ? mu_x2_addr1 : mu_x2_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35652_q <= 12'b000000000000;
    else
      n35652_q <= n35651_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n35653_o = instruction_tid_valid_in ? mu_y_addr1 : mu_y_addr1_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35654_q <= 12'b000000000000;
    else
      n35654_q <= n35653_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35655_q <= 1'b0;
    else
      n35655_q <= instruction_vm_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35656_q <= 1'b0;
    else
      n35656_q <= vm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35657_q <= 1'b0;
    else
      n35657_q <= vm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35658_q <= 1'b0;
    else
      n35658_q <= vm_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35659_q <= 1'b0;
    else
      n35659_q <= vm_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35660_q <= 1'b0;
    else
      n35660_q <= vm_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35662_q <= 5'b00000;
    else
      n35662_q <= imu_opcode;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35663_q <= 4'b0000;
    else
      n35663_q <= imu_x1_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35664_q <= 4'b0000;
    else
      n35664_q <= imu_x2_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35665_q <= 4'b0000;
    else
      n35665_q <= imu_y_parm;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35666_q <= 13'b0000000000000;
    else
      n35666_q <= imu_const;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35667_q <= 5'b00000;
    else
      n35667_q <= imu_opcode_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35668_q <= 4'b0000;
    else
      n35668_q <= imu_x1_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35669_q <= 4'b0000;
    else
      n35669_q <= imu_x2_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35670_q <= 4'b0000;
    else
      n35670_q <= imu_y_parm_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35671_q <= 4'b0000;
    else
      n35671_q <= imu_x1_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35672_q <= 4'b0000;
    else
      n35672_q <= imu_x2_parm_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35673_q <= 13'b0000000000000;
    else
      n35673_q <= imu_const_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35674_q <= 13'b0000000000000;
    else
      n35674_q <= imu_const_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35675_q <= 3'b000;
    else
      n35675_q <= n34933_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35676_q <= 3'b000;
    else
      n35676_q <= imu_y_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35677_q <= 3'b000;
    else
      n35677_q <= imu_y_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35678_q <= 3'b000;
    else
      n35678_q <= imu_y_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35680_q <= 1'b0;
    else
      n35680_q <= n34935_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35681_q <= 1'b0;
    else
      n35681_q <= imu_y_valid_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35682_q <= 1'b0;
    else
      n35682_q <= imu_y_valid_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35683_q <= 1'b0;
    else
      n35683_q <= imu_y_valid_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35685_q <= 5'b00000;
    else
      n35685_q <= n34937_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  always @(posedge clock_in or posedge n34841_o)
    if (n34841_o)
      n35686_q <= 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n35686_q <= n34865_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35687_q <= 13'b0000000000000;
    else
      n35687_q <= n35764_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35688_q <= 13'b0000000000000;
    else
      n35688_q <= n35778_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35689_q <= 13'b0000000000000;
    else
      n35689_q <= imu_x1_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35690_q <= 13'b0000000000000;
    else
      n35690_q <= imu_x2_ireg_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35691_q <= 13'b0000000000000;
    else
      n35691_q <= imu_x1_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35692_q <= 13'b0000000000000;
    else
      n35692_q <= imu_x2_ireg_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35693_q <= 8'b00000000;
    else
      n35693_q <= n35544_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35694_q <= 8'b00000000;
    else
      n35694_q <= mu_lane_r;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35695_q <= 8'b00000000;
    else
      n35695_q <= mu_lane_rr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35696_q <= 8'b00000000;
    else
      n35696_q <= mu_lane_rrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35697_q <= 8'b00000000;
    else
      n35697_q <= mu_lane_rrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35698_q <= 8'b00000000;
    else
      n35698_q <= mu_lane_rrrrr;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35699_q <= 8'b00000000;
    else
      n35699_q <= n35546_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35700_q <= 8'b00000000;
    else
      n35700_q <= n35548_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  always @(posedge clock_in or posedge n35516_o)
    if (n35516_o)
      n35701_q <= 8'b00000000;
    else
      n35701_q <= n35550_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  always @(posedge clock_in or posedge n34898_o)
    if (n34898_o)
      n35702_q <= 13'b0000000000000;
    else
      n35702_q <= result_in;
  /* ../../HW/src/pcore/instr_decoder2.vhd:114:16  */
  assign n35703_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:113:16  */
  assign n35704_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:109:16  */
  assign n35705_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:108:16  */
  assign n35706_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n35707_o = n34772_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  always @*
    case (n35707_o)
      2'b00: n35708_o = n35703_o;
      2'b01: n35708_o = n35704_o;
      2'b10: n35708_o = n35705_o;
      2'b11: n35708_o = n35706_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:28  */
  assign n35709_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:455:29  */
  assign n35710_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:100:16  */
  assign n35711_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:99:16  */
  assign n35712_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n35713_o = n34782_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  always @*
    case (n35713_o)
      2'b00: n35714_o = n35709_o;
      2'b01: n35714_o = n35710_o;
      2'b10: n35714_o = n35711_o;
      2'b11: n35714_o = n35712_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:28  */
  assign n35715_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:456:29  */
  assign n35716_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:96:16  */
  assign n35717_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:94:16  */
  assign n35718_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n35719_o = n34792_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  always @*
    case (n35719_o)
      2'b00: n35720_o = n35715_o;
      2'b01: n35720_o = n35716_o;
      2'b10: n35720_o = n35717_o;
      2'b11: n35720_o = n35718_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:28  */
  assign n35721_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:457:29  */
  assign n35722_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:89:16  */
  assign n35723_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:88:16  */
  assign n35724_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n35725_o = n34802_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  always @*
    case (n35725_o)
      2'b00: n35726_o = n35721_o;
      2'b01: n35726_o = n35722_o;
      2'b10: n35726_o = n35723_o;
      2'b11: n35726_o = n35724_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:28  */
  assign n35727_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:459:29  */
  assign n35728_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:82:16  */
  assign n35729_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:81:16  */
  assign n35730_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n35731_o = n34806_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  always @*
    case (n35731_o)
      2'b00: n35732_o = n35727_o;
      2'b01: n35732_o = n35728_o;
      2'b10: n35732_o = n35729_o;
      2'b11: n35732_o = n35730_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:28  */
  assign n35733_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:460:29  */
  assign n35734_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:76:16  */
  assign n35735_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:73:16  */
  assign n35736_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n35737_o = n34811_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  always @*
    case (n35737_o)
      2'b00: n35738_o = n35733_o;
      2'b01: n35738_o = n35734_o;
      2'b10: n35738_o = n35735_o;
      2'b11: n35738_o = n35736_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:28  */
  assign n35739_o = iregisters_lo[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:463:29  */
  assign n35740_o = iregisters_lo[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:69:16  */
  assign n35741_o = iregisters_lo[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:66:16  */
  assign n35742_o = iregisters_lo[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n35743_o = n34819_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  always @*
    case (n35743_o)
      2'b00: n35744_o = n35739_o;
      2'b01: n35744_o = n35740_o;
      2'b10: n35744_o = n35741_o;
      2'b11: n35744_o = n35742_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:27  */
  assign n35745_o = iregisters_hi[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:466:28  */
  assign n35746_o = iregisters_hi[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n35747_o = iregisters_hi[38:26];
  /* ../../HW/src/pcore/instr_decoder2.vhd:609:5  */
  assign n35748_o = iregisters_hi[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n35749_o = n34829_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  always @*
    case (n35749_o)
      2'b00: n35750_o = n35745_o;
      2'b01: n35750_o = n35746_o;
      2'b10: n35750_o = n35747_o;
      2'b11: n35750_o = n35748_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:27  */
  assign n35751_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:467:28  */
  assign n35752_o = iregisters_r[25:13];
  /* ../../HW/src/pcore/instr_decoder2.vhd:510:5  */
  assign n35753_o = iregisters_r[38:26];
  assign n35754_o = iregisters_r[51:39];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n35755_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n35756_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:738:9  */
  assign n35757_o = iregisters_r[90:78];
  /* ../../HW/src/pcore/instr_decoder2.vhd:711:1  */
  assign n35758_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n35759_o = n34900_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n35759_o)
      2'b00: n35760_o = n35751_o;
      2'b01: n35760_o = n35752_o;
      2'b10: n35760_o = n35753_o;
      2'b11: n35760_o = n35754_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n35761_o = n34900_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  always @*
    case (n35761_o)
      2'b00: n35762_o = n35755_o;
      2'b01: n35762_o = n35756_o;
      2'b10: n35762_o = n35757_o;
      2'b11: n35762_o = n35758_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n35763_o = n34900_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n35764_o = n35763_o ? n35762_o : n35760_o;
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:38  */
  assign n35765_o = iregisters_r[12:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:619:39  */
  assign n35766_o = iregisters_r[25:13];
  assign n35767_o = iregisters_r[38:26];
  assign n35768_o = iregisters_r[51:39];
  assign n35769_o = iregisters_r[64:52];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:50  */
  assign n35770_o = iregisters_r[77:65];
  /* ../../HW/src/pcore/instr_decoder2.vhd:308:60  */
  assign n35771_o = iregisters_r[90:78];
  assign n35772_o = iregisters_r[103:91];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n35773_o = n34904_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n35773_o)
      2'b00: n35774_o = n35765_o;
      2'b01: n35774_o = n35766_o;
      2'b10: n35774_o = n35767_o;
      2'b11: n35774_o = n35768_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n35775_o = n34904_o[1:0];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  always @*
    case (n35775_o)
      2'b00: n35776_o = n35769_o;
      2'b01: n35776_o = n35770_o;
      2'b10: n35776_o = n35771_o;
      2'b11: n35776_o = n35772_o;
    endcase
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n35777_o = n34904_o[2];
  /* ../../HW/src/pcore/instr_decoder2.vhd:620:38  */
  assign n35778_o = n35777_o ? n35776_o : n35774_o;
endmodule

module register_bank
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  rd_en_in,
   input  rd_en_vm_in,
   input  rd_x1_vector_in,
   input  [11:0] rd_x1_addr_in,
   input  rd_x2_vector_in,
   input  [11:0] rd_x2_addr_in,
   input  wr_en_in,
   input  wr_en_vm_in,
   input  wr_vector_in,
   input  [11:0] wr_addr_in,
   input  [95:0] wr_data_in,
   input  [7:0] wr_lane_in,
   input  [2:0] dp_rd_vector_in,
   input  [1:0] dp_rd_scatter_in,
   input  [2:0] dp_rd_scatter_cnt_in,
   input  [2:0] dp_rd_scatter_vector_in,
   input  dp_rd_gen_valid_in,
   input  [1:0] dp_rd_data_flow_in,
   input  [1:0] dp_rd_data_type_in,
   input  dp_rd_stream_in,
   input  [1:0] dp_rd_stream_id_in,
   input  [16:0] dp_rd_addr_in,
   input  [2:0] dp_wr_vector_in,
   input  [16:0] dp_wr_addr_in,
   input  dp_write_in,
   input  dp_write_vm_in,
   input  dp_read_in,
   input  dp_read_vm_in,
   input  [95:0] dp_writedata_in,
   output rd_en_out,
   output [95:0] rd_x1_data_out,
   output [95:0] rd_x2_data_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output [1:0] dp_read_scatter_out,
   output [2:0] dp_read_scatter_cnt_out,
   output [2:0] dp_read_scatter_vector_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire rd_en_vm1;
  wire rd_en_vm2;
  wire wr_en_vm1;
  wire wr_en_vm2;
  wire dp_read_vm1;
  wire dp_read_vm2;
  wire dp_write_vm1;
  wire dp_write_vm2;
  wire dp_readena_vm1;
  wire dp_readena_vm2;
  wire [11:0] dp_encode;
  wire [95:0] dp_readdata_vm;
  wire [95:0] dp_readdata_vm1;
  wire [95:0] dp_readdata_vm2;
  wire [11:0] q1_encode;
  wire [11:0] q2_encode;
  wire [95:0] rd_x1_data_vm;
  wire [95:0] rd_x2_data_vm;
  wire [95:0] rd_x1_data1_vm1;
  wire [95:0] rd_x2_data1_vm1;
  wire [95:0] rd_x1_data1_vm2;
  wire [95:0] rd_x2_data1_vm2;
  wire rd_enable1_vm1;
  wire rd_enable1_vm2;
  wire [1:0] dp_rd_data_flow_r;
  wire [1:0] dp_rd_data_type_r;
  wire dp_rd_stream_r;
  wire [1:0] dp_rd_stream_id_r;
  wire dp_rd_gen_valid_r;
  wire [1:0] dp_rd_scatter_r;
  wire [2:0] dp_rd_scatter_cnt_r;
  wire [2:0] dp_rd_scatter_vector_r;
  wire [2:0] dp_rd_vaddr_r;
  wire [2:0] dp_rd_vector_r;
  wire [1:0] dp_rd_data_flow_rr;
  wire [1:0] dp_rd_data_type_rr;
  wire dp_rd_stream_rr;
  wire [1:0] dp_rd_stream_id_rr;
  wire dp_rd_gen_valid_rr;
  wire [1:0] dp_rd_scatter_rr;
  wire [2:0] dp_rd_scatter_cnt_rr;
  wire [2:0] dp_rd_scatter_vector_rr;
  wire [2:0] dp_rd_vaddr_rr;
  wire [2:0] dp_rd_vector_rr;
  wire rd_x1_vector_r;
  wire rd_x1_vector_rr;
  wire [2:0] rd_x1_vaddr_r;
  wire [2:0] rd_x1_vaddr_rr;
  wire rd_x2_vector_r;
  wire rd_x2_vector_rr;
  wire [2:0] rd_x2_vaddr_r;
  wire [2:0] rd_x2_vaddr_rr;
  wire n34326_o;
  wire n34327_o;
  wire n34328_o;
  wire n34329_o;
  wire n34330_o;
  wire n34331_o;
  wire n34332_o;
  wire n34333_o;
  wire n34334_o;
  wire n34335_o;
  wire n34336_o;
  wire n34337_o;
  wire [83:0] n34338_o;
  wire n34340_o;
  wire n34342_o;
  wire n34346_o;
  wire [23:0] n34347_o;
  wire [35:0] n34348_o;
  wire [47:0] n34349_o;
  wire [59:0] n34350_o;
  wire [71:0] n34351_o;
  wire [83:0] n34352_o;
  wire [95:0] n34353_o;
  wire [95:0] n34354_o;
  wire n34356_o;
  wire [23:0] n34357_o;
  wire [35:0] n34358_o;
  wire [47:0] n34359_o;
  wire [59:0] n34360_o;
  wire [71:0] n34361_o;
  wire [83:0] n34362_o;
  wire [95:0] n34363_o;
  wire [95:0] n34364_o;
  wire n34366_o;
  wire n34369_o;
  wire [2:0] n34372_o;
  wire [2:0] n34373_o;
  wire [2:0] n34374_o;
  wire [95:0] n34460_o;
  wire [11:0] n34464_o;
  wire n34466_o;
  wire [11:0] n34467_o;
  wire n34469_o;
  wire [11:0] n34470_o;
  wire n34472_o;
  wire [11:0] n34473_o;
  wire n34475_o;
  wire [11:0] n34476_o;
  wire n34478_o;
  wire [11:0] n34479_o;
  wire n34481_o;
  wire [11:0] n34482_o;
  wire n34484_o;
  wire [11:0] n34485_o;
  wire [6:0] n34486_o;
  reg [11:0] n34487_o;
  wire [95:0] n34489_o;
  wire [11:0] n34493_o;
  wire n34495_o;
  wire [11:0] n34496_o;
  wire n34498_o;
  wire [11:0] n34499_o;
  wire n34501_o;
  wire [11:0] n34502_o;
  wire n34504_o;
  wire [11:0] n34505_o;
  wire n34507_o;
  wire [11:0] n34508_o;
  wire n34510_o;
  wire [11:0] n34511_o;
  wire n34513_o;
  wire [11:0] n34514_o;
  wire [6:0] n34515_o;
  reg [11:0] n34516_o;
  wire [95:0] n34518_o;
  wire [11:0] n34522_o;
  wire n34524_o;
  wire [11:0] n34525_o;
  wire n34527_o;
  wire [11:0] n34528_o;
  wire n34530_o;
  wire [11:0] n34531_o;
  wire n34533_o;
  wire [11:0] n34534_o;
  wire n34536_o;
  wire [11:0] n34537_o;
  wire n34539_o;
  wire [11:0] n34540_o;
  wire n34542_o;
  wire [11:0] n34543_o;
  wire [6:0] n34544_o;
  reg [11:0] n34545_o;
  wire register_file_i_n34547;
  wire [95:0] register_file_i_n34548;
  wire [95:0] register_file_i_n34549;
  wire [95:0] register_file_i_n34550;
  wire register_file_i_n34551;
  wire register_file_i_rd_en_out;
  wire [95:0] register_file_i_rd_x1_data_out;
  wire [95:0] register_file_i_rd_x2_data_out;
  wire [95:0] register_file_i_dp_readdata_out;
  wire register_file_i_dp_readena_out;
  wire register_file_i2_n34562;
  wire [95:0] register_file_i2_n34563;
  wire [95:0] register_file_i2_n34564;
  wire [95:0] register_file_i2_n34565;
  wire register_file_i2_n34566;
  wire register_file_i2_rd_en_out;
  wire [95:0] register_file_i2_rd_x1_data_out;
  wire [95:0] register_file_i2_rd_x2_data_out;
  wire [95:0] register_file_i2_dp_readdata_out;
  wire register_file_i2_dp_readena_out;
  reg [1:0] n34599_q;
  reg [1:0] n34600_q;
  reg n34601_q;
  reg [1:0] n34602_q;
  reg n34603_q;
  reg [1:0] n34604_q;
  reg [2:0] n34605_q;
  reg [2:0] n34606_q;
  reg [2:0] n34607_q;
  reg [2:0] n34608_q;
  reg [1:0] n34609_q;
  reg [1:0] n34610_q;
  reg n34611_q;
  reg [1:0] n34612_q;
  reg n34613_q;
  reg [1:0] n34614_q;
  reg [2:0] n34615_q;
  reg [2:0] n34616_q;
  reg [2:0] n34617_q;
  reg [2:0] n34618_q;
  reg n34619_q;
  reg n34620_q;
  reg [2:0] n34621_q;
  reg [2:0] n34622_q;
  reg n34623_q;
  reg n34624_q;
  reg [2:0] n34625_q;
  reg [2:0] n34626_q;
  wire [95:0] n34627_o;
  assign rd_en_out = n34342_o;
  assign rd_x1_data_out = n34354_o;
  assign rd_x2_data_out = n34364_o;
  assign dp_readdata_out = n34627_o;
  assign dp_readdata_vm_out = n34340_o;
  assign dp_readena_out = n34366_o;
  assign dp_read_vector_out = dp_rd_vector_rr;
  assign dp_read_vaddr_out = dp_rd_vaddr_rr;
  assign dp_read_scatter_out = dp_rd_scatter_rr;
  assign dp_read_scatter_cnt_out = dp_rd_scatter_cnt_rr;
  assign dp_read_scatter_vector_out = dp_rd_scatter_vector_rr;
  assign dp_read_gen_valid_out = dp_rd_gen_valid_rr;
  assign dp_read_data_flow_out = dp_rd_data_flow_rr;
  assign dp_read_data_type_out = dp_rd_data_type_rr;
  assign dp_read_stream_out = dp_rd_stream_rr;
  assign dp_read_stream_id_out = dp_rd_stream_id_rr;
  /* ../../HW/src/pcore/register_bank.vhd:117:8  */
  assign rd_en_vm1 = n34327_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:118:8  */
  assign rd_en_vm2 = n34328_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:119:8  */
  assign wr_en_vm1 = n34330_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:120:8  */
  assign wr_en_vm2 = n34331_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:121:8  */
  assign dp_read_vm1 = n34333_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:122:8  */
  assign dp_read_vm2 = n34334_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:123:8  */
  assign dp_write_vm1 = n34336_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:124:8  */
  assign dp_write_vm2 = n34337_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:125:8  */
  assign dp_readena_vm1 = register_file_i_n34551; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:126:8  */
  assign dp_readena_vm2 = register_file_i2_n34566; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:141:8  */
  assign dp_encode = n34487_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:144:8  */
  assign dp_readdata_vm = n34460_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:145:8  */
  assign dp_readdata_vm1 = register_file_i_n34550; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:146:8  */
  assign dp_readdata_vm2 = register_file_i2_n34565; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:147:8  */
  assign q1_encode = n34516_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:148:8  */
  assign q2_encode = n34545_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:149:8  */
  assign rd_x1_data_vm = n34489_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:150:8  */
  assign rd_x2_data_vm = n34518_o; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:151:8  */
  assign rd_x1_data1_vm1 = register_file_i_n34548; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:152:8  */
  assign rd_x2_data1_vm1 = register_file_i_n34549; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:153:8  */
  assign rd_x1_data1_vm2 = register_file_i2_n34563; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:154:8  */
  assign rd_x2_data1_vm2 = register_file_i2_n34564; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:155:8  */
  assign rd_enable1_vm1 = register_file_i_n34547; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:156:8  */
  assign rd_enable1_vm2 = register_file_i2_n34562; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:164:8  */
  assign dp_rd_data_flow_r = n34599_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:165:8  */
  assign dp_rd_data_type_r = n34600_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:166:8  */
  assign dp_rd_stream_r = n34601_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:167:8  */
  assign dp_rd_stream_id_r = n34602_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:168:8  */
  assign dp_rd_gen_valid_r = n34603_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:169:8  */
  assign dp_rd_scatter_r = n34604_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:170:8  */
  assign dp_rd_scatter_cnt_r = n34605_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:171:8  */
  assign dp_rd_scatter_vector_r = n34606_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:172:8  */
  assign dp_rd_vaddr_r = n34607_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:173:8  */
  assign dp_rd_vector_r = n34608_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:175:8  */
  assign dp_rd_data_flow_rr = n34609_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:176:8  */
  assign dp_rd_data_type_rr = n34610_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:177:8  */
  assign dp_rd_stream_rr = n34611_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:178:8  */
  assign dp_rd_stream_id_rr = n34612_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:179:8  */
  assign dp_rd_gen_valid_rr = n34613_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:180:8  */
  assign dp_rd_scatter_rr = n34614_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:181:8  */
  assign dp_rd_scatter_cnt_rr = n34615_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:182:8  */
  assign dp_rd_scatter_vector_rr = n34616_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:183:8  */
  assign dp_rd_vaddr_rr = n34617_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:184:8  */
  assign dp_rd_vector_rr = n34618_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:186:8  */
  assign rd_x1_vector_r = n34619_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:187:8  */
  assign rd_x1_vector_rr = n34620_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:188:8  */
  assign rd_x1_vaddr_r = n34621_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:189:8  */
  assign rd_x1_vaddr_rr = n34622_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:190:8  */
  assign rd_x2_vector_r = n34623_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:191:8  */
  assign rd_x2_vector_rr = n34624_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:192:8  */
  assign rd_x2_vaddr_r = n34625_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:193:8  */
  assign rd_x2_vaddr_rr = n34626_q; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:197:28  */
  assign n34326_o = ~rd_en_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:197:23  */
  assign n34327_o = rd_en_in & n34326_o;
  /* ../../HW/src/pcore/register_bank.vhd:198:23  */
  assign n34328_o = rd_en_in & rd_en_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:200:28  */
  assign n34329_o = ~wr_en_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:200:23  */
  assign n34330_o = wr_en_in & n34329_o;
  /* ../../HW/src/pcore/register_bank.vhd:201:23  */
  assign n34331_o = wr_en_in & wr_en_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:203:32  */
  assign n34332_o = ~dp_read_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:203:27  */
  assign n34333_o = dp_read_in & n34332_o;
  /* ../../HW/src/pcore/register_bank.vhd:204:27  */
  assign n34334_o = dp_read_in & dp_read_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:205:34  */
  assign n34335_o = ~dp_write_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:205:29  */
  assign n34336_o = dp_write_in & n34335_o;
  /* ../../HW/src/pcore/register_bank.vhd:206:29  */
  assign n34337_o = dp_write_in & dp_write_vm_in;
  /* ../../HW/src/pcore/register_bank.vhd:209:84  */
  assign n34338_o = dp_readdata_vm[95:12];
  /* ../../HW/src/pcore/register_bank.vhd:211:27  */
  assign n34340_o = dp_readena_vm1 ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/register_bank.vhd:213:29  */
  assign n34342_o = rd_enable1_vm1 | rd_enable1_vm2;
  /* ../../HW/src/pcore/register_bank.vhd:221:22  */
  assign n34346_o = rd_x1_vector_rr != 1'b0;
  /* ../../HW/src/pcore/register_bank.vhd:224:35  */
  assign n34347_o = {q1_encode, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:225:35  */
  assign n34348_o = {n34347_o, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:226:35  */
  assign n34349_o = {n34348_o, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:227:35  */
  assign n34350_o = {n34349_o, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:228:35  */
  assign n34351_o = {n34350_o, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:229:35  */
  assign n34352_o = {n34351_o, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:230:35  */
  assign n34353_o = {n34352_o, q1_encode};
  /* ../../HW/src/pcore/register_bank.vhd:221:4  */
  assign n34354_o = n34346_o ? rd_x1_data_vm : n34353_o;
  /* ../../HW/src/pcore/register_bank.vhd:233:22  */
  assign n34356_o = rd_x2_vector_rr != 1'b0;
  /* ../../HW/src/pcore/register_bank.vhd:236:35  */
  assign n34357_o = {q2_encode, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:237:35  */
  assign n34358_o = {n34357_o, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:238:35  */
  assign n34359_o = {n34358_o, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:239:35  */
  assign n34360_o = {n34359_o, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:240:35  */
  assign n34361_o = {n34360_o, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:241:35  */
  assign n34362_o = {n34361_o, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:242:35  */
  assign n34363_o = {n34362_o, q2_encode};
  /* ../../HW/src/pcore/register_bank.vhd:233:4  */
  assign n34364_o = n34356_o ? rd_x2_data_vm : n34363_o;
  /* ../../HW/src/pcore/register_bank.vhd:247:34  */
  assign n34366_o = dp_readena_vm1 | dp_readena_vm2;
  /* ../../HW/src/pcore/register_bank.vhd:261:17  */
  assign n34369_o = ~reset_in;
  /* ../../HW/src/pcore/register_bank.vhd:320:41  */
  assign n34372_o = rd_x1_addr_in[2:0];
  /* ../../HW/src/pcore/register_bank.vhd:324:41  */
  assign n34373_o = rd_x2_addr_in[2:0];
  /* ../../HW/src/pcore/register_bank.vhd:327:41  */
  assign n34374_o = dp_rd_addr_in[2:0];
  /* ../../HW/src/pcore/register_bank.vhd:332:36  */
  assign n34460_o = dp_readena_vm1 ? dp_readdata_vm1 : dp_readdata_vm2;
  /* ../../HW/src/pcore/register_bank.vhd:343:34  */
  assign n34464_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/register_bank.vhd:342:4  */
  assign n34466_o = dp_rd_vaddr_rr == 3'b000;
  /* ../../HW/src/pcore/register_bank.vhd:345:34  */
  assign n34467_o = dp_readdata_vm[23:12];
  /* ../../HW/src/pcore/register_bank.vhd:344:4  */
  assign n34469_o = dp_rd_vaddr_rr == 3'b001;
  /* ../../HW/src/pcore/register_bank.vhd:347:34  */
  assign n34470_o = dp_readdata_vm[35:24];
  /* ../../HW/src/pcore/register_bank.vhd:346:4  */
  assign n34472_o = dp_rd_vaddr_rr == 3'b010;
  /* ../../HW/src/pcore/register_bank.vhd:349:34  */
  assign n34473_o = dp_readdata_vm[47:36];
  /* ../../HW/src/pcore/register_bank.vhd:348:4  */
  assign n34475_o = dp_rd_vaddr_rr == 3'b011;
  /* ../../HW/src/pcore/register_bank.vhd:351:34  */
  assign n34476_o = dp_readdata_vm[59:48];
  /* ../../HW/src/pcore/register_bank.vhd:350:4  */
  assign n34478_o = dp_rd_vaddr_rr == 3'b100;
  /* ../../HW/src/pcore/register_bank.vhd:353:34  */
  assign n34479_o = dp_readdata_vm[71:60];
  /* ../../HW/src/pcore/register_bank.vhd:352:4  */
  assign n34481_o = dp_rd_vaddr_rr == 3'b101;
  /* ../../HW/src/pcore/register_bank.vhd:355:34  */
  assign n34482_o = dp_readdata_vm[83:72];
  /* ../../HW/src/pcore/register_bank.vhd:354:4  */
  assign n34484_o = dp_rd_vaddr_rr == 3'b110;
  /* ../../HW/src/pcore/register_bank.vhd:357:34  */
  assign n34485_o = dp_readdata_vm[95:84];
  assign n34486_o = {n34484_o, n34481_o, n34478_o, n34475_o, n34472_o, n34469_o, n34466_o};
  /* ../../HW/src/pcore/register_bank.vhd:341:1  */
  always @*
    case (n34486_o)
      7'b1000000: n34487_o = n34482_o;
      7'b0100000: n34487_o = n34479_o;
      7'b0010000: n34487_o = n34476_o;
      7'b0001000: n34487_o = n34473_o;
      7'b0000100: n34487_o = n34470_o;
      7'b0000010: n34487_o = n34467_o;
      7'b0000001: n34487_o = n34464_o;
      default: n34487_o = n34485_o;
    endcase
  /* ../../HW/src/pcore/register_bank.vhd:362:34  */
  assign n34489_o = rd_enable1_vm1 ? rd_x1_data1_vm1 : rd_x1_data1_vm2;
  /* ../../HW/src/pcore/register_bank.vhd:373:33  */
  assign n34493_o = rd_x1_data_vm[11:0];
  /* ../../HW/src/pcore/register_bank.vhd:372:4  */
  assign n34495_o = rd_x1_vaddr_rr == 3'b000;
  /* ../../HW/src/pcore/register_bank.vhd:375:33  */
  assign n34496_o = rd_x1_data_vm[23:12];
  /* ../../HW/src/pcore/register_bank.vhd:374:4  */
  assign n34498_o = rd_x1_vaddr_rr == 3'b001;
  /* ../../HW/src/pcore/register_bank.vhd:377:33  */
  assign n34499_o = rd_x1_data_vm[35:24];
  /* ../../HW/src/pcore/register_bank.vhd:376:4  */
  assign n34501_o = rd_x1_vaddr_rr == 3'b010;
  /* ../../HW/src/pcore/register_bank.vhd:379:33  */
  assign n34502_o = rd_x1_data_vm[47:36];
  /* ../../HW/src/pcore/register_bank.vhd:378:4  */
  assign n34504_o = rd_x1_vaddr_rr == 3'b011;
  /* ../../HW/src/pcore/register_bank.vhd:381:33  */
  assign n34505_o = rd_x1_data_vm[59:48];
  /* ../../HW/src/pcore/register_bank.vhd:380:4  */
  assign n34507_o = rd_x1_vaddr_rr == 3'b100;
  /* ../../HW/src/pcore/register_bank.vhd:383:33  */
  assign n34508_o = rd_x1_data_vm[71:60];
  /* ../../HW/src/pcore/register_bank.vhd:382:4  */
  assign n34510_o = rd_x1_vaddr_rr == 3'b101;
  /* ../../HW/src/pcore/register_bank.vhd:385:33  */
  assign n34511_o = rd_x1_data_vm[83:72];
  /* ../../HW/src/pcore/register_bank.vhd:384:4  */
  assign n34513_o = rd_x1_vaddr_rr == 3'b110;
  /* ../../HW/src/pcore/register_bank.vhd:387:33  */
  assign n34514_o = rd_x1_data_vm[95:84];
  assign n34515_o = {n34513_o, n34510_o, n34507_o, n34504_o, n34501_o, n34498_o, n34495_o};
  /* ../../HW/src/pcore/register_bank.vhd:371:1  */
  always @*
    case (n34515_o)
      7'b1000000: n34516_o = n34511_o;
      7'b0100000: n34516_o = n34508_o;
      7'b0010000: n34516_o = n34505_o;
      7'b0001000: n34516_o = n34502_o;
      7'b0000100: n34516_o = n34499_o;
      7'b0000010: n34516_o = n34496_o;
      7'b0000001: n34516_o = n34493_o;
      default: n34516_o = n34514_o;
    endcase
  /* ../../HW/src/pcore/register_bank.vhd:392:34  */
  assign n34518_o = rd_enable1_vm1 ? rd_x2_data1_vm1 : rd_x2_data1_vm2;
  /* ../../HW/src/pcore/register_bank.vhd:403:33  */
  assign n34522_o = rd_x2_data_vm[11:0];
  /* ../../HW/src/pcore/register_bank.vhd:402:4  */
  assign n34524_o = rd_x2_vaddr_rr == 3'b000;
  /* ../../HW/src/pcore/register_bank.vhd:405:33  */
  assign n34525_o = rd_x2_data_vm[23:12];
  /* ../../HW/src/pcore/register_bank.vhd:404:4  */
  assign n34527_o = rd_x2_vaddr_rr == 3'b001;
  /* ../../HW/src/pcore/register_bank.vhd:407:33  */
  assign n34528_o = rd_x2_data_vm[35:24];
  /* ../../HW/src/pcore/register_bank.vhd:406:4  */
  assign n34530_o = rd_x2_vaddr_rr == 3'b010;
  /* ../../HW/src/pcore/register_bank.vhd:409:33  */
  assign n34531_o = rd_x2_data_vm[47:36];
  /* ../../HW/src/pcore/register_bank.vhd:408:4  */
  assign n34533_o = rd_x2_vaddr_rr == 3'b011;
  /* ../../HW/src/pcore/register_bank.vhd:411:33  */
  assign n34534_o = rd_x2_data_vm[59:48];
  /* ../../HW/src/pcore/register_bank.vhd:410:4  */
  assign n34536_o = rd_x2_vaddr_rr == 3'b100;
  /* ../../HW/src/pcore/register_bank.vhd:413:33  */
  assign n34537_o = rd_x2_data_vm[71:60];
  /* ../../HW/src/pcore/register_bank.vhd:412:4  */
  assign n34539_o = rd_x2_vaddr_rr == 3'b101;
  /* ../../HW/src/pcore/register_bank.vhd:415:33  */
  assign n34540_o = rd_x2_data_vm[83:72];
  /* ../../HW/src/pcore/register_bank.vhd:414:4  */
  assign n34542_o = rd_x2_vaddr_rr == 3'b110;
  /* ../../HW/src/pcore/register_bank.vhd:417:33  */
  assign n34543_o = rd_x2_data_vm[95:84];
  assign n34544_o = {n34542_o, n34539_o, n34536_o, n34533_o, n34530_o, n34527_o, n34524_o};
  /* ../../HW/src/pcore/register_bank.vhd:401:1  */
  always @*
    case (n34544_o)
      7'b1000000: n34545_o = n34540_o;
      7'b0100000: n34545_o = n34537_o;
      7'b0010000: n34545_o = n34534_o;
      7'b0001000: n34545_o = n34531_o;
      7'b0000100: n34545_o = n34528_o;
      7'b0000010: n34545_o = n34525_o;
      7'b0000001: n34545_o = n34522_o;
      default: n34545_o = n34543_o;
    endcase
  /* ../../HW/src/pcore/register_bank.vhd:431:46  */
  assign register_file_i_n34547 = register_file_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:436:50  */
  assign register_file_i_n34548 = register_file_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:437:50  */
  assign register_file_i_n34549 = register_file_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:461:52  */
  assign register_file_i_n34550 = register_file_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:462:51  */
  assign register_file_i_n34551 = register_file_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:425:1  */
  register_file register_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en_vm1),
    .rd_x1_vector_in(rd_x1_vector_in),
    .rd_x1_addr_in(rd_x1_addr_in),
    .rd_x2_vector_in(rd_x2_vector_in),
    .rd_x2_addr_in(rd_x2_addr_in),
    .wr_en_in(wr_en_vm1),
    .wr_vector_in(wr_vector_in),
    .wr_addr_in(wr_addr_in),
    .wr_data_in(wr_data_in),
    .wr_lane_in(wr_lane_in),
    .dp_rd_vector_in(dp_rd_vector_in),
    .dp_rd_scatter_in(dp_rd_scatter_in),
    .dp_rd_scatter_cnt_in(dp_rd_scatter_cnt_in),
    .dp_rd_scatter_vector_in(dp_rd_scatter_vector_in),
    .dp_rd_gen_valid_in(dp_rd_gen_valid_in),
    .dp_rd_data_flow_in(dp_rd_data_flow_in),
    .dp_rd_data_type_in(dp_rd_data_type_in),
    .dp_rd_stream_in(dp_rd_stream_in),
    .dp_rd_stream_id_in(dp_rd_stream_id_in),
    .dp_rd_addr_in(dp_rd_addr_in),
    .dp_wr_vector_in(dp_wr_vector_in),
    .dp_wr_addr_in(dp_wr_addr_in),
    .dp_write_in(dp_write_vm1),
    .dp_read_in(dp_read_vm1),
    .dp_writedata_in(dp_writedata_in),
    .rd_en_out(register_file_i_rd_en_out),
    .rd_x1_data_out(register_file_i_rd_x1_data_out),
    .rd_x2_data_out(register_file_i_rd_x2_data_out),
    .dp_readdata_out(register_file_i_dp_readdata_out),
    .dp_readena_out(register_file_i_dp_readena_out));
  /* ../../HW/src/pcore/register_bank.vhd:475:46  */
  assign register_file_i2_n34562 = register_file_i2_rd_en_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:480:50  */
  assign register_file_i2_n34563 = register_file_i2_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:481:50  */
  assign register_file_i2_n34564 = register_file_i2_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:505:52  */
  assign register_file_i2_n34565 = register_file_i2_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:506:51  */
  assign register_file_i2_n34566 = register_file_i2_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/register_bank.vhd:469:1  */
  register_file register_file_i2 (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en_vm2),
    .rd_x1_vector_in(rd_x1_vector_in),
    .rd_x1_addr_in(rd_x1_addr_in),
    .rd_x2_vector_in(rd_x2_vector_in),
    .rd_x2_addr_in(rd_x2_addr_in),
    .wr_en_in(wr_en_vm2),
    .wr_vector_in(wr_vector_in),
    .wr_addr_in(wr_addr_in),
    .wr_data_in(wr_data_in),
    .wr_lane_in(wr_lane_in),
    .dp_rd_vector_in(dp_rd_vector_in),
    .dp_rd_scatter_in(dp_rd_scatter_in),
    .dp_rd_scatter_cnt_in(dp_rd_scatter_cnt_in),
    .dp_rd_scatter_vector_in(dp_rd_scatter_vector_in),
    .dp_rd_gen_valid_in(dp_rd_gen_valid_in),
    .dp_rd_data_flow_in(dp_rd_data_flow_in),
    .dp_rd_data_type_in(dp_rd_data_type_in),
    .dp_rd_stream_in(dp_rd_stream_in),
    .dp_rd_stream_id_in(dp_rd_stream_id_in),
    .dp_rd_addr_in(dp_rd_addr_in),
    .dp_wr_vector_in(dp_wr_vector_in),
    .dp_wr_addr_in(dp_wr_addr_in),
    .dp_write_in(dp_write_vm2),
    .dp_read_in(dp_read_vm2),
    .dp_writedata_in(dp_writedata_in),
    .rd_en_out(register_file_i2_rd_en_out),
    .rd_x1_data_out(register_file_i2_rd_x1_data_out),
    .rd_x2_data_out(register_file_i2_rd_x2_data_out),
    .dp_readdata_out(register_file_i2_dp_readdata_out),
    .dp_readena_out(register_file_i2_dp_readena_out));
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34599_q <= 2'b00;
    else
      n34599_q <= dp_rd_data_flow_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34600_q <= 2'b00;
    else
      n34600_q <= dp_rd_data_type_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34601_q <= 1'b0;
    else
      n34601_q <= dp_rd_stream_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34602_q <= 2'b00;
    else
      n34602_q <= dp_rd_stream_id_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34603_q <= 1'b0;
    else
      n34603_q <= dp_rd_gen_valid_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34604_q <= 2'b00;
    else
      n34604_q <= dp_rd_scatter_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34605_q <= 3'b000;
    else
      n34605_q <= dp_rd_scatter_cnt_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34606_q <= 3'b000;
    else
      n34606_q <= dp_rd_scatter_vector_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34607_q <= 3'b000;
    else
      n34607_q <= n34374_o;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34608_q <= 3'b000;
    else
      n34608_q <= dp_rd_vector_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34609_q <= 2'b00;
    else
      n34609_q <= dp_rd_data_flow_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34610_q <= 2'b00;
    else
      n34610_q <= dp_rd_data_type_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34611_q <= 1'b0;
    else
      n34611_q <= dp_rd_stream_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34612_q <= 2'b00;
    else
      n34612_q <= dp_rd_stream_id_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34613_q <= 1'b0;
    else
      n34613_q <= dp_rd_gen_valid_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34614_q <= 2'b00;
    else
      n34614_q <= dp_rd_scatter_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34615_q <= 3'b000;
    else
      n34615_q <= dp_rd_scatter_cnt_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34616_q <= 3'b000;
    else
      n34616_q <= dp_rd_scatter_vector_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34617_q <= 3'b000;
    else
      n34617_q <= dp_rd_vaddr_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34618_q <= 3'b000;
    else
      n34618_q <= dp_rd_vector_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34619_q <= 1'b0;
    else
      n34619_q <= rd_x1_vector_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34620_q <= 1'b0;
    else
      n34620_q <= rd_x1_vector_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34621_q <= 3'b000;
    else
      n34621_q <= n34372_o;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34622_q <= 3'b000;
    else
      n34622_q <= rd_x1_vaddr_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34623_q <= 1'b0;
    else
      n34623_q <= rd_x2_vector_in;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34624_q <= 1'b0;
    else
      n34624_q <= rd_x2_vector_r;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34625_q <= 3'b000;
    else
      n34625_q <= n34373_o;
  /* ../../HW/src/pcore/register_bank.vhd:295:8  */
  always @(posedge clock_in or posedge n34369_o)
    if (n34369_o)
      n34626_q <= 3'b000;
    else
      n34626_q <= rd_x2_vaddr_r;
  /* ../../HW/src/pcore/register_bank.vhd:261:5  */
  assign n34627_o = {n34338_o, dp_encode};
endmodule

module ialu
  (input  clock_in,
   input  reset_in,
   input  [4:0] opcode_in,
   input  [12:0] x1_in,
   input  [12:0] x2_in,
   output [12:0] y_out,
   output y_neg_out,
   output y_zero_out);
  wire [12:0] x1;
  wire [12:0] x2;
  wire [12:0] shift_y;
  wire [12:0] logic_shift_y;
  wire [12:0] y_r;
  wire [12:0] y2_r;
  wire [12:0] x1_r;
  wire [12:0] x2_r;
  wire [4:0] opcode_r;
  wire [4:0] opcode_rr;
  wire [25:0] mul_y;
  wire [12:0] mul_x1;
  wire [12:0] mul_x2;
  wire shr;
  wire n34223_o;
  wire n34224_o;
  wire [25:0] mult_i_n34226;
  wire [25:0] mult_i_z_out;
  wire [3:0] n34229_o;
  wire [12:0] shifter_i_n34230;
  wire [12:0] shifter_i_data_out;
  localparam n34233_o = 1'b1;
  wire [3:0] n34234_o;
  wire [12:0] logic_shifter_i_n34235;
  wire [12:0] logic_shifter_i_data_out;
  wire n34238_o;
  wire n34241_o;
  wire n34242_o;
  wire n34246_o;
  wire [12:0] n34248_o;
  wire n34250_o;
  wire [12:0] n34251_o;
  wire n34253_o;
  wire n34255_o;
  wire n34257_o;
  wire n34258_o;
  wire n34260_o;
  wire [12:0] n34261_o;
  wire n34263_o;
  wire [12:0] n34264_o;
  wire n34266_o;
  wire [12:0] n34267_o;
  wire n34269_o;
  wire [6:0] n34270_o;
  reg [12:0] n34272_o;
  wire [12:0] n34273_o;
  wire n34275_o;
  reg [12:0] n34276_o;
  reg [12:0] n34302_q;
  reg [12:0] n34303_q;
  reg [12:0] n34305_q;
  reg [12:0] n34306_q;
  reg [4:0] n34307_q;
  reg [4:0] n34308_q;
  assign y_out = y_r;
  assign y_neg_out = n34238_o;
  assign y_zero_out = n34242_o;
  /* ../../HW/src/ialu/ialu.vhd:45:8  */
  assign x1 = x1_r; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:46:8  */
  assign x2 = x2_r; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:47:8  */
  assign shift_y = shifter_i_n34230; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:48:8  */
  assign logic_shift_y = logic_shifter_i_n34235; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:49:8  */
  assign y_r = n34302_q; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:50:8  */
  assign y2_r = n34303_q; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:52:8  */
  assign x1_r = n34305_q; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:53:8  */
  assign x2_r = n34306_q; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:54:8  */
  assign opcode_r = n34307_q; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:55:8  */
  assign opcode_rr = n34308_q; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:57:8  */
  assign mul_y = mult_i_n34226; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:58:8  */
  assign mul_x1 = x1_r; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:59:8  */
  assign mul_x2 = x2_r; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:60:8  */
  assign shr = n34224_o; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:69:26  */
  assign n34223_o = opcode_r == 5'b00100;
  /* ../../HW/src/ialu/ialu.vhd:69:12  */
  assign n34224_o = n34223_o ? 1'b0 : 1'b1;
  /* ../../HW/src/ialu/ialu.vhd:87:16  */
  assign mult_i_n34226 = mult_i_z_out; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:75:1  */
  multiplier_13_bf8b4530d8d246dd74ac53a13471bba17941dff7 mult_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .x_in(mul_x1),
    .y_in(mul_x2),
    .z_out(mult_i_z_out));
  /* ../../HW/src/ialu/ialu.vhd:102:22  */
  assign n34229_o = x2[3:0];
  /* ../../HW/src/ialu/ialu.vhd:103:17  */
  assign shifter_i_n34230 = shifter_i_data_out; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:94:1  */
  barrel_shifter_a_4_13 shifter_i (
    .direction_in(shr),
    .data_in(x1),
    .distance_in(n34229_o),
    .data_out(shifter_i_data_out));
  /* ../../HW/src/ialu/ialu.vhd:114:22  */
  assign n34234_o = x2[3:0];
  /* ../../HW/src/ialu/ialu.vhd:115:17  */
  assign logic_shifter_i_n34235 = logic_shifter_i_data_out; // (signal)
  /* ../../HW/src/ialu/ialu.vhd:106:1  */
  barrel_shifter_l_4_13 logic_shifter_i (
    .direction_in(n34233_o),
    .data_in(x1),
    .distance_in(n34234_o),
    .data_out(logic_shifter_i_data_out));
  /* ../../HW/src/ialu/ialu.vhd:119:17  */
  assign n34238_o = y_r[12];
  /* ../../HW/src/ialu/ialu.vhd:120:27  */
  assign n34241_o = y_r == 13'b0000000000000;
  /* ../../HW/src/ialu/ialu.vhd:120:19  */
  assign n34242_o = n34241_o ? 1'b1 : 1'b0;
  /* ../../HW/src/ialu/ialu.vhd:124:12  */
  assign n34246_o = ~reset_in;
  /* ../../HW/src/ialu/ialu.vhd:149:29  */
  assign n34248_o = x1_r + x2_r;
  /* ../../HW/src/ialu/ialu.vhd:148:13  */
  assign n34250_o = opcode_r == 5'b00001;
  /* ../../HW/src/ialu/ialu.vhd:151:29  */
  assign n34251_o = x1_r - x2_r;
  /* ../../HW/src/ialu/ialu.vhd:150:13  */
  assign n34253_o = opcode_r == 5'b00010;
  /* ../../HW/src/ialu/ialu.vhd:152:13  */
  assign n34255_o = opcode_r == 5'b00100;
  /* ../../HW/src/ialu/ialu.vhd:152:34  */
  assign n34257_o = opcode_r == 5'b00101;
  /* ../../HW/src/ialu/ialu.vhd:152:34  */
  assign n34258_o = n34255_o | n34257_o;
  /* ../../HW/src/ialu/ialu.vhd:154:13  */
  assign n34260_o = opcode_r == 5'b01001;
  /* ../../HW/src/ialu/ialu.vhd:157:57  */
  assign n34261_o = x1_r | x2_r;
  /* ../../HW/src/ialu/ialu.vhd:156:13  */
  assign n34263_o = opcode_r == 5'b00110;
  /* ../../HW/src/ialu/ialu.vhd:159:57  */
  assign n34264_o = x1_r & x2_r;
  /* ../../HW/src/ialu/ialu.vhd:158:13  */
  assign n34266_o = opcode_r == 5'b00111;
  /* ../../HW/src/ialu/ialu.vhd:161:57  */
  assign n34267_o = x1_r ^ x2_r;
  /* ../../HW/src/ialu/ialu.vhd:160:13  */
  assign n34269_o = opcode_r == 5'b01000;
  /* ../../HW/src/alu/alu.vhd:306:5  */
  assign n34270_o = {n34269_o, n34266_o, n34263_o, n34260_o, n34258_o, n34253_o, n34250_o};
  /* ../../HW/src/ialu/ialu.vhd:147:9  */
  always @*
    case (n34270_o)
      7'b1000000: n34272_o = n34267_o;
      7'b0100000: n34272_o = n34264_o;
      7'b0010000: n34272_o = n34261_o;
      7'b0001000: n34272_o = logic_shift_y;
      7'b0000100: n34272_o = shift_y;
      7'b0000010: n34272_o = n34251_o;
      7'b0000001: n34272_o = n34248_o;
      default: n34272_o = 13'b0000000000000;
    endcase
  /* ../../HW/src/ialu/ialu.vhd:172:38  */
  assign n34273_o = mul_y[12:0];
  /* ../../HW/src/ialu/ialu.vhd:171:13  */
  assign n34275_o = opcode_rr == 5'b00011;
  /* ../../HW/src/ialu/ialu.vhd:170:9  */
  always @*
    case (n34275_o)
      1'b1: n34276_o = n34273_o;
      default: n34276_o = y2_r;
    endcase
  /* ../../HW/src/ialu/ialu.vhd:134:5  */
  always @(posedge clock_in or posedge n34246_o)
    if (n34246_o)
      n34302_q <= 13'b0000000000000;
    else
      n34302_q <= n34276_o;
  /* ../../HW/src/ialu/ialu.vhd:134:5  */
  always @(posedge clock_in or posedge n34246_o)
    if (n34246_o)
      n34303_q <= 13'b0000000000000;
    else
      n34303_q <= n34272_o;
  /* ../../HW/src/ialu/ialu.vhd:134:5  */
  always @(posedge clock_in or posedge n34246_o)
    if (n34246_o)
      n34305_q <= 13'b0000000000000;
    else
      n34305_q <= x1_in;
  /* ../../HW/src/ialu/ialu.vhd:134:5  */
  always @(posedge clock_in or posedge n34246_o)
    if (n34246_o)
      n34306_q <= 13'b0000000000000;
    else
      n34306_q <= x2_in;
  /* ../../HW/src/ialu/ialu.vhd:134:5  */
  always @(posedge clock_in or posedge n34246_o)
    if (n34246_o)
      n34307_q <= 5'b00000;
    else
      n34307_q <= opcode_in;
  /* ../../HW/src/ialu/ialu.vhd:134:5  */
  always @(posedge clock_in or posedge n34246_o)
    if (n34246_o)
      n34308_q <= 5'b00000;
    else
      n34308_q <= opcode_r;
endmodule

module alu
  (input  clock_in,
   input  reset_in,
   input  [4:0] mu_opcode_in,
   input  [3:0] mu_tid_in,
   input  [31:0] xreg_in,
   input  [11:0] x1_in,
   input  [11:0] x2_in,
   input  [11:0] x_scalar_in,
   output [31:0] y_out,
   output y2_out,
   output [11:0] y3_out);
  wire add_sub_r;
  wire [31:0] y_add;
  wire [31:0] y_add_r;
  wire [23:0] y_mul;
  wire negative;
  wire zero;
  wire [31:0] y_r;
  wire y2_r;
  wire [11:0] y3_r;
  wire [31:0] xreg_r;
  wire [31:0] xreg_rr;
  wire [4:0] mu_opcode_r;
  wire [4:0] mu_opcode_rr;
  wire [4:0] mu_opcode_rrr;
  wire [4:0] mu_opcode_rrrr;
  wire [11:0] mul_x2_r;
  wire [11:0] x1_r;
  wire [11:0] x2_r;
  wire [11:0] x_scalar_r;
  wire [31:0] y_shift;
  wire [31:0] y_shift_r;
  wire [1:0] shift_distance_r;
  wire [1:0] shift_distance_rr;
  wire shift_direction_r;
  wire shift_direction_rr;
  wire [7:0] y_mul_ext;
  wire [31:0] add_x1;
  wire n33833_o;
  wire n33836_o;
  wire n33837_o;
  wire n33841_o;
  wire n33843_o;
  wire n33844_o;
  wire n33846_o;
  wire n33847_o;
  wire n33849_o;
  wire n33850_o;
  wire n33851_o;
  wire n33852_o;
  wire n33854_o;
  wire n33855_o;
  wire n33856_o;
  wire n33858_o;
  wire n33860_o;
  wire n33861_o;
  wire n33863_o;
  wire n33864_o;
  wire [5:0] n33865_o;
  reg n33866_o;
  wire [8:0] n33867_o;
  wire n33869_o;
  wire [8:0] n33870_o;
  wire n33872_o;
  wire [31:0] n33874_o;
  wire [31:0] n33876_o;
  wire n33883_o;
  wire n33884_o;
  wire [20:0] n33885_o;
  wire n33887_o;
  wire [11:0] n33888_o;
  wire [11:0] n33890_o;
  wire [20:0] n33891_o;
  wire n33893_o;
  wire [11:0] n33894_o;
  wire [11:0] n33896_o;
  wire [11:0] n33897_o;
  wire [23:0] mul_i_n33909;
  wire [23:0] mul_i_z_out;
  wire [31:0] adder_i_n33912;
  wire [31:0] adder_i_z_out;
  wire [31:0] shifter_i_n33915;
  wire [31:0] shifter_i_data_out;
  wire n33918_o;
  wire n33919_o;
  wire n33920_o;
  wire n33921_o;
  wire n33922_o;
  wire n33923_o;
  wire n33924_o;
  wire n33925_o;
  wire [3:0] n33926_o;
  wire [3:0] n33927_o;
  wire [7:0] n33928_o;
  wire [31:0] n33929_o;
  wire n33932_o;
  wire n33935_o;
  wire [1:0] n33936_o;
  wire n33938_o;
  wire n33940_o;
  wire n33942_o;
  wire n33943_o;
  wire n33945_o;
  wire n33946_o;
  wire n33948_o;
  wire n33949_o;
  wire [11:0] n33952_o;
  wire [11:0] n33953_o;
  wire [11:0] n33954_o;
  wire n33961_o;
  wire n33964_o;
  wire n33966_o;
  wire n33967_o;
  wire n33969_o;
  wire n33970_o;
  wire n33972_o;
  wire n33973_o;
  wire n33974_o;
  wire [9:0] n33975_o;
  wire n33977_o;
  wire [1:0] n33978_o;
  wire [1:0] n33980_o;
  wire [1:0] n33982_o;
  wire [1:0] n33984_o;
  wire n33986_o;
  wire n33988_o;
  wire n33989_o;
  wire n33992_o;
  wire n34020_o;
  wire [1:0] n34022_o;
  wire n34024_o;
  wire n34026_o;
  wire n34028_o;
  wire n34029_o;
  wire n34031_o;
  wire n34033_o;
  wire n34034_o;
  wire n34036_o;
  wire n34037_o;
  wire n34038_o;
  wire n34039_o;
  wire n34040_o;
  wire n34041_o;
  wire n34042_o;
  wire n34043_o;
  wire n34044_o;
  wire n34045_o;
  wire n34046_o;
  wire n34047_o;
  wire n34048_o;
  wire n34049_o;
  wire n34050_o;
  wire n34051_o;
  wire n34052_o;
  wire n34053_o;
  wire n34054_o;
  wire n34055_o;
  wire n34056_o;
  wire n34057_o;
  wire [3:0] n34058_o;
  wire [3:0] n34059_o;
  wire [3:0] n34060_o;
  wire [3:0] n34061_o;
  wire [3:0] n34062_o;
  wire [15:0] n34063_o;
  wire [19:0] n34064_o;
  wire n34066_o;
  wire n34068_o;
  wire n34069_o;
  wire n34070_o;
  wire n34071_o;
  wire n34072_o;
  wire n34073_o;
  wire n34074_o;
  wire n34075_o;
  wire n34076_o;
  wire n34077_o;
  wire n34078_o;
  wire n34079_o;
  wire n34080_o;
  wire n34081_o;
  wire n34082_o;
  wire n34083_o;
  wire n34084_o;
  wire n34085_o;
  wire n34086_o;
  wire n34087_o;
  wire n34088_o;
  wire n34089_o;
  wire [3:0] n34090_o;
  wire [3:0] n34091_o;
  wire [3:0] n34092_o;
  wire [3:0] n34093_o;
  wire [3:0] n34094_o;
  wire [15:0] n34095_o;
  wire [19:0] n34096_o;
  wire [2:0] n34097_o;
  wire [11:0] n34098_o;
  reg [11:0] n34100_o;
  wire [19:0] n34101_o;
  reg [19:0] n34103_o;
  wire [31:0] n34104_o;
  wire [31:0] n34105_o;
  wire [1:0] n34106_o;
  wire n34108_o;
  wire n34109_o;
  wire n34110_o;
  wire n34112_o;
  wire n34114_o;
  wire n34116_o;
  wire n34118_o;
  wire n34119_o;
  wire n34121_o;
  wire n34122_o;
  wire n34124_o;
  wire n34125_o;
  wire n34127_o;
  wire n34128_o;
  wire n34130_o;
  wire n34131_o;
  wire [2:0] n34132_o;
  reg n34137_o;
  wire n34138_o;
  reg n34189_q;
  reg [31:0] n34190_q;
  reg [31:0] n34191_q;
  reg n34192_q;
  reg [11:0] n34193_q;
  reg [31:0] n34194_q;
  reg [31:0] n34195_q;
  reg [4:0] n34198_q;
  reg [4:0] n34199_q;
  reg [4:0] n34200_q;
  reg [4:0] n34201_q;
  reg [11:0] n34204_q;
  reg [11:0] n34205_q;
  reg [11:0] n34206_q;
  reg [11:0] n34207_q;
  reg [31:0] n34208_q;
  reg [1:0] n34210_q;
  reg [1:0] n34211_q;
  reg n34214_q;
  reg n34215_q;
  assign y_out = y_r;
  assign y2_out = y2_r;
  assign y3_out = y3_r;
  /* ../../HW/src/alu/alu.vhd:51:8  */
  assign add_sub_r = n34189_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:52:8  */
  assign y_add = adder_i_n33912; // (signal)
  /* ../../HW/src/alu/alu.vhd:53:8  */
  assign y_add_r = n34190_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:54:8  */
  assign y_mul = mul_i_n33909; // (signal)
  /* ../../HW/src/alu/alu.vhd:55:8  */
  assign negative = n33833_o; // (signal)
  /* ../../HW/src/alu/alu.vhd:56:8  */
  assign zero = n33837_o; // (signal)
  /* ../../HW/src/alu/alu.vhd:57:8  */
  assign y_r = n34191_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:58:8  */
  assign y2_r = n34192_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:59:8  */
  assign y3_r = n34193_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:63:8  */
  assign xreg_r = n34194_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:64:8  */
  assign xreg_rr = n34195_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:70:8  */
  assign mu_opcode_r = n34198_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:71:8  */
  assign mu_opcode_rr = n34199_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:72:8  */
  assign mu_opcode_rrr = n34200_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:73:8  */
  assign mu_opcode_rrrr = n34201_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:77:8  */
  assign mul_x2_r = n34204_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:78:8  */
  assign x1_r = n34205_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:79:8  */
  assign x2_r = n34206_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:80:8  */
  assign x_scalar_r = n34207_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:88:8  */
  assign y_shift = shifter_i_n33915; // (signal)
  /* ../../HW/src/alu/alu.vhd:89:8  */
  assign y_shift_r = n34208_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:91:8  */
  assign shift_distance_r = n34210_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:92:8  */
  assign shift_distance_rr = n34211_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:95:8  */
  assign shift_direction_r = n34214_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:96:8  */
  assign shift_direction_rr = n34215_q; // (signal)
  /* ../../HW/src/alu/alu.vhd:99:8  */
  assign y_mul_ext = n33928_o; // (signal)
  /* ../../HW/src/alu/alu.vhd:100:8  */
  assign add_x1 = n33929_o; // (signal)
  /* ../../HW/src/alu/alu.vhd:137:22  */
  assign n33833_o = y_shift_r[31];
  /* ../../HW/src/alu/alu.vhd:139:27  */
  assign n33836_o = y_shift_r == 32'b00000000000000000000000000000000;
  /* ../../HW/src/alu/alu.vhd:139:13  */
  assign n33837_o = n33836_o ? 1'b1 : 1'b0;
  /* ../../HW/src/alu/alu.vhd:153:16  */
  assign n33841_o = ~reset_in;
  /* ../../HW/src/alu/alu.vhd:161:33  */
  assign n33843_o = ~zero;
  /* ../../HW/src/alu/alu.vhd:161:28  */
  assign n33844_o = negative & n33843_o;
  /* ../../HW/src/alu/alu.vhd:160:7  */
  assign n33846_o = mu_opcode_rrrr == 5'b00110;
  /* ../../HW/src/alu/alu.vhd:163:28  */
  assign n33847_o = negative | zero;
  /* ../../HW/src/alu/alu.vhd:162:7  */
  assign n33849_o = mu_opcode_rrrr == 5'b00111;
  /* ../../HW/src/alu/alu.vhd:165:20  */
  assign n33850_o = ~negative;
  /* ../../HW/src/alu/alu.vhd:165:39  */
  assign n33851_o = ~zero;
  /* ../../HW/src/alu/alu.vhd:165:34  */
  assign n33852_o = n33850_o & n33851_o;
  /* ../../HW/src/alu/alu.vhd:164:7  */
  assign n33854_o = mu_opcode_rrrr == 5'b01000;
  /* ../../HW/src/alu/alu.vhd:167:20  */
  assign n33855_o = ~negative;
  /* ../../HW/src/alu/alu.vhd:167:34  */
  assign n33856_o = n33855_o | zero;
  /* ../../HW/src/alu/alu.vhd:166:7  */
  assign n33858_o = mu_opcode_rrrr == 5'b01001;
  /* ../../HW/src/alu/alu.vhd:168:7  */
  assign n33860_o = mu_opcode_rrrr == 5'b01010;
  /* ../../HW/src/alu/alu.vhd:171:18  */
  assign n33861_o = ~zero;
  /* ../../HW/src/alu/alu.vhd:170:7  */
  assign n33863_o = mu_opcode_rrrr == 5'b01011;
  /* ../../HW/src/alu/alu.vhd:173:27  */
  assign n33864_o = y_shift_r[0];
  assign n33865_o = {n33863_o, n33860_o, n33858_o, n33854_o, n33849_o, n33846_o};
  /* ../../HW/src/alu/alu.vhd:159:4  */
  always @*
    case (n33865_o)
      6'b100000: n33866_o = n33861_o;
      6'b010000: n33866_o = zero;
      6'b001000: n33866_o = n33856_o;
      6'b000100: n33866_o = n33852_o;
      6'b000010: n33866_o = n33847_o;
      6'b000001: n33866_o = n33844_o;
      default: n33866_o = n33864_o;
    endcase
  /* ../../HW/src/alu/alu.vhd:176:16  */
  assign n33867_o = y_shift_r[31:23];
  /* ../../HW/src/alu/alu.vhd:176:30  */
  assign n33869_o = n33867_o == 9'b011111111;
  /* ../../HW/src/alu/alu.vhd:179:19  */
  assign n33870_o = y_shift_r[31:23];
  /* ../../HW/src/alu/alu.vhd:179:33  */
  assign n33872_o = n33870_o == 9'b100000000;
  /* ../../HW/src/alu/alu.vhd:179:4  */
  assign n33874_o = n33872_o ? 32'b10000000100000000000000000000000 : y_shift_r;
  /* ../../HW/src/alu/alu.vhd:176:4  */
  assign n33876_o = n33869_o ? 32'b01111111100000000000000000000000 : n33874_o;
  /* ../../HW/src/alu/alu.vhd:114:15  */
  assign n33883_o = y_shift_r[31];
  /* ../../HW/src/alu/alu.vhd:114:38  */
  assign n33884_o = ~n33883_o;
  /* ../../HW/src/alu/alu.vhd:116:18  */
  assign n33885_o = y_shift_r[31:11];
  /* ../../HW/src/alu/alu.vhd:116:67  */
  assign n33887_o = n33885_o == 21'b000000000000000000000;
  /* ../../HW/src/alu/alu.vhd:117:30  */
  assign n33888_o = y_shift_r[11:0];
  /* ../../HW/src/alu/alu.vhd:116:7  */
  assign n33890_o = n33887_o ? n33888_o : 12'b011111111111;
  /* ../../HW/src/alu/alu.vhd:122:18  */
  assign n33891_o = y_shift_r[31:11];
  /* ../../HW/src/alu/alu.vhd:122:67  */
  assign n33893_o = n33891_o == 21'b111111111111111111111;
  /* ../../HW/src/alu/alu.vhd:123:30  */
  assign n33894_o = y_shift_r[11:0];
  /* ../../HW/src/alu/alu.vhd:122:7  */
  assign n33896_o = n33893_o ? n33894_o : 12'b100000000000;
  /* ../../HW/src/alu/alu.vhd:114:4  */
  assign n33897_o = n33884_o ? n33890_o : n33896_o;
  /* ../../HW/src/alu/alu.vhd:204:16  */
  assign mul_i_n33909 = mul_i_z_out; // (signal)
  /* ../../HW/src/alu/alu.vhd:192:1  */
  multiplier_12_bf8b4530d8d246dd74ac53a13471bba17941dff7 mul_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .x_in(x2_r),
    .y_in(mul_x2_r),
    .z_out(mul_i_z_out));
  /* ../../HW/src/alu/alu.vhd:217:14  */
  assign adder_i_n33912 = adder_i_z_out; // (signal)
  /* ../../HW/src/alu/alu.vhd:207:1  */
  adder_32 adder_i (
    .x_in(xreg_rr),
    .y_in(add_x1),
    .add_sub_in(add_sub_r),
    .z_out(adder_i_z_out));
  /* ../../HW/src/alu/alu.vhd:233:17  */
  assign shifter_i_n33915 = shifter_i_data_out; // (signal)
  /* ../../HW/src/alu/alu.vhd:224:1  */
  barrel_shifter_a_2_32 shifter_i (
    .direction_in(shift_direction_rr),
    .data_in(y_add_r),
    .distance_in(shift_distance_rr),
    .data_out(shifter_i_data_out));
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33918_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33919_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33920_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33921_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33922_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33923_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33924_o = y_mul[23];
  /* ../../HW/src/alu/alu.vhd:236:28  */
  assign n33925_o = y_mul[23];
  assign n33926_o = {n33918_o, n33919_o, n33920_o, n33921_o};
  assign n33927_o = {n33922_o, n33923_o, n33924_o, n33925_o};
  assign n33928_o = {n33926_o, n33927_o};
  /* ../../HW/src/alu/alu.vhd:238:21  */
  assign n33929_o = {y_mul_ext, y_mul};
  /* ../../HW/src/alu/alu.vhd:242:16  */
  assign n33932_o = ~reset_in;
  /* ../../HW/src/alu/alu.vhd:246:22  */
  assign n33935_o = mu_opcode_in == 5'b01100;
  /* ../../HW/src/alu/alu.vhd:248:25  */
  assign n33936_o = mu_opcode_in[4:3];
  /* ../../HW/src/alu/alu.vhd:248:55  */
  assign n33938_o = n33936_o == 2'b11;
  /* ../../HW/src/alu/alu.vhd:250:25  */
  assign n33940_o = mu_opcode_in == 5'b00010;
  /* ../../HW/src/alu/alu.vhd:251:22  */
  assign n33942_o = mu_opcode_in == 5'b00001;
  /* ../../HW/src/alu/alu.vhd:250:49  */
  assign n33943_o = n33940_o | n33942_o;
  /* ../../HW/src/alu/alu.vhd:252:22  */
  assign n33945_o = mu_opcode_in == 5'b10100;
  /* ../../HW/src/alu/alu.vhd:251:42  */
  assign n33946_o = n33943_o | n33945_o;
  /* ../../HW/src/alu/alu.vhd:253:22  */
  assign n33948_o = mu_opcode_in == 5'b10110;
  /* ../../HW/src/alu/alu.vhd:252:40  */
  assign n33949_o = n33946_o | n33948_o;
  /* ../../HW/src/alu/alu.vhd:250:7  */
  assign n33952_o = n33949_o ? 12'b000000000000 : 12'b000000000001;
  /* ../../HW/src/alu/alu.vhd:248:7  */
  assign n33953_o = n33938_o ? x1_in : n33952_o;
  /* ../../HW/src/alu/alu.vhd:246:7  */
  assign n33954_o = n33935_o ? x1_in : n33953_o;
  /* ../../HW/src/alu/alu.vhd:265:13  */
  assign n33961_o = ~reset_in;
  /* ../../HW/src/alu/alu.vhd:276:18  */
  assign n33964_o = mu_opcode_r == 5'b10110;
  /* ../../HW/src/alu/alu.vhd:276:50  */
  assign n33966_o = mu_opcode_r == 5'b10100;
  /* ../../HW/src/alu/alu.vhd:276:36  */
  assign n33967_o = n33964_o | n33966_o;
  /* ../../HW/src/alu/alu.vhd:276:82  */
  assign n33969_o = mu_opcode_r == 5'b10101;
  /* ../../HW/src/alu/alu.vhd:276:68  */
  assign n33970_o = n33967_o | n33969_o;
  /* ../../HW/src/alu/alu.vhd:276:113  */
  assign n33972_o = mu_opcode_r == 5'b10011;
  /* ../../HW/src/alu/alu.vhd:276:99  */
  assign n33973_o = n33970_o | n33972_o;
  /* ../../HW/src/alu/alu.vhd:278:20  */
  assign n33974_o = x_scalar_r[11];
  /* ../../HW/src/alu/alu.vhd:280:32  */
  assign n33975_o = x_scalar_r[11:2];
  /* ../../HW/src/alu/alu.vhd:280:82  */
  assign n33977_o = n33975_o != 10'b0000000000;
  /* ../../HW/src/alu/alu.vhd:283:40  */
  assign n33978_o = x_scalar_r[1:0];
  /* ../../HW/src/alu/alu.vhd:280:7  */
  assign n33980_o = n33977_o ? 2'b11 : n33978_o;
  /* ../../HW/src/alu/alu.vhd:278:7  */
  assign n33982_o = n33974_o ? 2'b00 : n33980_o;
  /* ../../HW/src/alu/alu.vhd:276:4  */
  assign n33984_o = n33973_o ? n33982_o : 2'b00;
  /* ../../HW/src/alu/alu.vhd:288:18  */
  assign n33986_o = mu_opcode_r == 5'b10100;
  /* ../../HW/src/alu/alu.vhd:288:50  */
  assign n33988_o = mu_opcode_r == 5'b10011;
  /* ../../HW/src/alu/alu.vhd:288:36  */
  assign n33989_o = n33986_o | n33988_o;
  /* ../../HW/src/alu/alu.vhd:288:4  */
  assign n33992_o = n33989_o ? 1'b0 : 1'b1;
  /* ../../HW/src/alu/alu.vhd:306:17  */
  assign n34020_o = ~reset_in;
  /* ../../HW/src/alu/alu.vhd:347:27  */
  assign n34022_o = mu_opcode_r[4:3];
  /* ../../HW/src/alu/alu.vhd:347:57  */
  assign n34024_o = n34022_o == 2'b11;
  /* ../../HW/src/alu/alu.vhd:351:19  */
  assign n34026_o = mu_opcode_r == 5'b10100;
  /* ../../HW/src/alu/alu.vhd:351:40  */
  assign n34028_o = mu_opcode_r == 5'b10110;
  /* ../../HW/src/alu/alu.vhd:351:40  */
  assign n34029_o = n34026_o | n34028_o;
  /* ../../HW/src/alu/alu.vhd:353:19  */
  assign n34031_o = mu_opcode_r == 5'b01100;
  /* ../../HW/src/alu/alu.vhd:353:39  */
  assign n34033_o = mu_opcode_r == 5'b10011;
  /* ../../HW/src/alu/alu.vhd:353:39  */
  assign n34034_o = n34031_o | n34033_o;
  /* ../../HW/src/alu/alu.vhd:353:55  */
  assign n34036_o = mu_opcode_r == 5'b10101;
  /* ../../HW/src/alu/alu.vhd:353:55  */
  assign n34037_o = n34034_o | n34036_o;
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34038_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34039_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34040_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34041_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34042_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34043_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34044_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34045_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34046_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34047_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34048_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34049_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34050_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34051_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34052_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34053_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34054_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34055_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34056_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:357:93  */
  assign n34057_o = x1_r[11];
  assign n34058_o = {n34038_o, n34039_o, n34040_o, n34041_o};
  assign n34059_o = {n34042_o, n34043_o, n34044_o, n34045_o};
  assign n34060_o = {n34046_o, n34047_o, n34048_o, n34049_o};
  assign n34061_o = {n34050_o, n34051_o, n34052_o, n34053_o};
  assign n34062_o = {n34054_o, n34055_o, n34056_o, n34057_o};
  assign n34063_o = {n34058_o, n34059_o, n34060_o, n34061_o};
  assign n34064_o = {n34063_o, n34062_o};
  /* ../../HW/src/alu/alu.vhd:355:19  */
  assign n34066_o = mu_opcode_r == 5'b00010;
  /* ../../HW/src/alu/alu.vhd:355:46  */
  assign n34068_o = mu_opcode_r == 5'b00001;
  /* ../../HW/src/alu/alu.vhd:355:46  */
  assign n34069_o = n34066_o | n34068_o;
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34070_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34071_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34072_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34073_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34074_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34075_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34076_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34077_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34078_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34079_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34080_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34081_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34082_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34083_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34084_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34085_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34086_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34087_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34088_o = x1_r[11];
  /* ../../HW/src/alu/alu.vhd:360:93  */
  assign n34089_o = x1_r[11];
  assign n34090_o = {n34070_o, n34071_o, n34072_o, n34073_o};
  assign n34091_o = {n34074_o, n34075_o, n34076_o, n34077_o};
  assign n34092_o = {n34078_o, n34079_o, n34080_o, n34081_o};
  assign n34093_o = {n34082_o, n34083_o, n34084_o, n34085_o};
  assign n34094_o = {n34086_o, n34087_o, n34088_o, n34089_o};
  assign n34095_o = {n34090_o, n34091_o, n34092_o, n34093_o};
  assign n34096_o = {n34095_o, n34094_o};
  assign n34097_o = {n34069_o, n34037_o, n34029_o};
  assign n34098_o = xreg_r[11:0];
  /* ../../HW/src/alu/alu.vhd:350:16  */
  always @*
    case (n34097_o)
      3'b100: n34100_o = x1_r;
      3'b010: n34100_o = 12'b000000000000;
      3'b001: n34100_o = n34098_o;
      default: n34100_o = x1_r;
    endcase
  assign n34101_o = xreg_r[31:12];
  /* ../../HW/src/alu/alu.vhd:350:16  */
  always @*
    case (n34097_o)
      3'b100: n34103_o = n34064_o;
      3'b010: n34103_o = 20'b00000000000000000000;
      3'b001: n34103_o = n34101_o;
      default: n34103_o = n34096_o;
    endcase
  assign n34104_o = {n34103_o, n34100_o};
  /* ../../HW/src/alu/alu.vhd:347:13  */
  assign n34105_o = n34024_o ? xreg_r : n34104_o;
  /* ../../HW/src/alu/alu.vhd:364:27  */
  assign n34106_o = mu_opcode_r[4:3];
  /* ../../HW/src/alu/alu.vhd:364:57  */
  assign n34108_o = n34106_o == 2'b11;
  /* ../../HW/src/alu/alu.vhd:365:45  */
  assign n34109_o = mu_opcode_r[1];
  /* ../../HW/src/alu/alu.vhd:365:30  */
  assign n34110_o = ~n34109_o;
  /* ../../HW/src/alu/alu.vhd:368:21  */
  assign n34112_o = mu_opcode_r == 5'b00011;
  /* ../../HW/src/alu/alu.vhd:370:21  */
  assign n34114_o = mu_opcode_r == 5'b00100;
  /* ../../HW/src/alu/alu.vhd:372:21  */
  assign n34116_o = mu_opcode_r == 5'b00110;
  /* ../../HW/src/alu/alu.vhd:372:45  */
  assign n34118_o = mu_opcode_r == 5'b00111;
  /* ../../HW/src/alu/alu.vhd:372:45  */
  assign n34119_o = n34116_o | n34118_o;
  /* ../../HW/src/alu/alu.vhd:373:44  */
  assign n34121_o = mu_opcode_r == 5'b01000;
  /* ../../HW/src/alu/alu.vhd:373:44  */
  assign n34122_o = n34119_o | n34121_o;
  /* ../../HW/src/alu/alu.vhd:374:44  */
  assign n34124_o = mu_opcode_r == 5'b01001;
  /* ../../HW/src/alu/alu.vhd:374:44  */
  assign n34125_o = n34122_o | n34124_o;
  /* ../../HW/src/alu/alu.vhd:375:44  */
  assign n34127_o = mu_opcode_r == 5'b01010;
  /* ../../HW/src/alu/alu.vhd:375:44  */
  assign n34128_o = n34125_o | n34127_o;
  /* ../../HW/src/alu/alu.vhd:376:44  */
  assign n34130_o = mu_opcode_r == 5'b01011;
  /* ../../HW/src/alu/alu.vhd:376:44  */
  assign n34131_o = n34128_o | n34130_o;
  assign n34132_o = {n34131_o, n34114_o, n34112_o};
  /* ../../HW/src/alu/alu.vhd:367:17  */
  always @*
    case (n34132_o)
      3'b100: n34137_o = 1'b0;
      3'b010: n34137_o = 1'b0;
      3'b001: n34137_o = 1'b1;
      default: n34137_o = 1'b1;
    endcase
  /* ../../HW/src/alu/alu.vhd:364:13  */
  assign n34138_o = n34108_o ? n34110_o : n34137_o;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34189_q <= 1'b0;
    else
      n34189_q <= n34138_o;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34190_q <= 32'b00000000000000000000000000000000;
    else
      n34190_q <= y_add;
  /* ../../HW/src/alu/alu.vhd:158:4  */
  always @(posedge clock_in or posedge n33841_o)
    if (n33841_o)
      n34191_q <= 32'b00000000000000000000000000000000;
    else
      n34191_q <= n33876_o;
  /* ../../HW/src/alu/alu.vhd:158:4  */
  always @(posedge clock_in or posedge n33841_o)
    if (n33841_o)
      n34192_q <= 1'b0;
    else
      n34192_q <= n33866_o;
  /* ../../HW/src/alu/alu.vhd:158:4  */
  always @(posedge clock_in or posedge n33841_o)
    if (n33841_o)
      n34193_q <= 12'b000000000000;
    else
      n34193_q <= n33897_o;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34194_q <= 32'b00000000000000000000000000000000;
    else
      n34194_q <= xreg_in;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34195_q <= 32'b00000000000000000000000000000000;
    else
      n34195_q <= n34105_o;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34198_q <= 5'b00000;
    else
      n34198_q <= mu_opcode_in;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34199_q <= 5'b00000;
    else
      n34199_q <= mu_opcode_r;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34200_q <= 5'b00000;
    else
      n34200_q <= mu_opcode_rr;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34201_q <= 5'b00000;
    else
      n34201_q <= mu_opcode_rrr;
  /* ../../HW/src/alu/alu.vhd:245:4  */
  always @(posedge clock_in or posedge n33932_o)
    if (n33932_o)
      n34204_q <= 12'b000000000000;
    else
      n34204_q <= n33954_o;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34205_q <= 12'b000000000000;
    else
      n34205_q <= x1_in;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34206_q <= 12'b000000000000;
    else
      n34206_q <= x2_in;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34207_q <= 12'b000000000000;
    else
      n34207_q <= x_scalar_in;
  /* ../../HW/src/alu/alu.vhd:329:9  */
  always @(posedge clock_in or posedge n34020_o)
    if (n34020_o)
      n34208_q <= 32'b00000000000000000000000000000000;
    else
      n34208_q <= y_shift;
  /* ../../HW/src/alu/alu.vhd:275:4  */
  always @(posedge clock_in or posedge n33961_o)
    if (n33961_o)
      n34210_q <= 2'b00;
    else
      n34210_q <= n33984_o;
  /* ../../HW/src/alu/alu.vhd:275:4  */
  always @(posedge clock_in or posedge n33961_o)
    if (n33961_o)
      n34211_q <= 2'b00;
    else
      n34211_q <= shift_distance_r;
  /* ../../HW/src/alu/alu.vhd:275:4  */
  always @(posedge clock_in or posedge n33961_o)
    if (n33961_o)
      n34214_q <= 1'b0;
    else
      n34214_q <= n33992_o;
  /* ../../HW/src/alu/alu.vhd:275:4  */
  always @(posedge clock_in or posedge n33961_o)
    if (n33961_o)
      n34215_q <= 1'b0;
    else
      n34215_q <= shift_direction_r;
endmodule

module iregister_file
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  rd_en1_in,
   input  rd_vm_in,
   input  [3:0] rd_tid1_in,
   input  [3:0] wr_tid1_in,
   input  wr_en1_in,
   input  wr_vm_in,
   input  wr_lane_in,
   input  [2:0] wr_addr1_in,
   input  [12:0] wr_data1_in,
   output [103:0] rd_data1_out,
   output [12:0] rd_lane_out);
  wire [143:0] q1;
  wire [143:0] wrdata1;
  wire [17:0] byteena1;
  wire [4:0] rdaddr1;
  wire [4:0] wraddr1;
  wire [12:0] rd_lane_r;
  wire [4:0] n33729_o;
  wire [4:0] n33730_o;
  wire [12:0] n33733_o;
  wire [12:0] n33734_o;
  wire [12:0] n33735_o;
  wire [12:0] n33736_o;
  wire [12:0] n33737_o;
  wire [12:0] n33738_o;
  wire [12:0] n33739_o;
  wire [12:0] n33740_o;
  wire n33744_o;
  wire [12:0] n33746_o;
  wire [12:0] n33747_o;
  wire [30:0] n33754_o;
  wire [31:0] n33755_o;
  wire n33757_o;
  wire [1:0] n33758_o;
  wire [1:0] n33760_o;
  wire [30:0] n33761_o;
  wire [31:0] n33762_o;
  wire n33764_o;
  wire [1:0] n33765_o;
  wire [1:0] n33767_o;
  wire [30:0] n33768_o;
  wire [31:0] n33769_o;
  wire n33771_o;
  wire [1:0] n33772_o;
  wire [1:0] n33774_o;
  wire [30:0] n33775_o;
  wire [31:0] n33776_o;
  wire n33778_o;
  wire [1:0] n33779_o;
  wire [1:0] n33781_o;
  wire [30:0] n33782_o;
  wire [31:0] n33783_o;
  wire n33785_o;
  wire [1:0] n33786_o;
  wire [1:0] n33788_o;
  wire [30:0] n33789_o;
  wire [31:0] n33790_o;
  wire n33792_o;
  wire [1:0] n33793_o;
  wire [1:0] n33795_o;
  wire [30:0] n33796_o;
  wire [31:0] n33797_o;
  wire n33799_o;
  wire [1:0] n33800_o;
  wire [1:0] n33802_o;
  wire [30:0] n33803_o;
  wire [31:0] n33804_o;
  wire n33806_o;
  wire [1:0] n33807_o;
  wire [1:0] n33809_o;
  wire [12:0] n33810_o;
  wire [1:0] n33811_o;
  localparam n33813_o = 1'b1;
  wire [143:0] iregister_ram_i_n33814;
  wire [143:0] iregister_ram_i_q1_out;
  wire [143:0] n33826_o;
  wire [17:0] n33827_o;
  reg [12:0] n33828_q;
  wire [103:0] n33829_o;
  assign rd_data1_out = n33829_o;
  assign rd_lane_out = rd_lane_r;
  /* ../../HW/src/ialu/iregister_file.vhd:58:8  */
  assign q1 = iregister_ram_i_n33814; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:59:8  */
  assign wrdata1 = n33826_o; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:60:8  */
  assign byteena1 = n33827_o; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:61:8  */
  assign rdaddr1 = n33729_o; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:62:8  */
  assign wraddr1 = n33730_o; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:63:8  */
  assign rd_lane_r = n33828_q; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:101:21  */
  assign n33729_o = {rd_vm_in, rd_tid1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:102:21  */
  assign n33730_o = {wr_vm_in, wr_tid1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33733_o = q1[12:0];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33734_o = q1[28:16];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33735_o = q1[44:32];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33736_o = q1[60:48];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33737_o = q1[76:64];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33738_o = q1[92:80];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33739_o = q1[108:96];
  /* ../../HW/src/ialu/iregister_file.vhd:113:35  */
  assign n33740_o = q1[124:112];
  /* ../../HW/src/ialu/iregister_file.vhd:119:12  */
  assign n33744_o = ~reset_in;
  /* ../../HW/src/ialu/iregister_file.vhd:123:37  */
  assign n33746_o = q1[140:128];
  /* ../../HW/src/ialu/iregister_file.vhd:123:31  */
  assign n33747_o = ~n33746_o;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33754_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33755_o = {1'b0, n33754_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33757_o = 32'b00000000000000000000000000000000 == n33755_o;
  assign n33758_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33760_o = n33757_o ? n33758_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33761_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33762_o = {1'b0, n33761_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33764_o = 32'b00000000000000000000000000000001 == n33762_o;
  assign n33765_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33767_o = n33764_o ? n33765_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33768_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33769_o = {1'b0, n33768_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33771_o = 32'b00000000000000000000000000000010 == n33769_o;
  assign n33772_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33774_o = n33771_o ? n33772_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33775_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33776_o = {1'b0, n33775_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33778_o = 32'b00000000000000000000000000000011 == n33776_o;
  assign n33779_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33781_o = n33778_o ? n33779_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33782_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33783_o = {1'b0, n33782_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33785_o = 32'b00000000000000000000000000000100 == n33783_o;
  assign n33786_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33788_o = n33785_o ? n33786_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33789_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33790_o = {1'b0, n33789_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33792_o = 32'b00000000000000000000000000000101 == n33790_o;
  assign n33793_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33795_o = n33792_o ? n33793_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33796_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33797_o = {1'b0, n33796_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33799_o = 32'b00000000000000000000000000000110 == n33797_o;
  assign n33800_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33802_o = n33799_o ? n33800_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:137:10  */
  assign n33803_o = {28'b0, wr_addr1_in};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33804_o = {1'b0, n33803_o};  //  uext
  /* ../../HW/src/ialu/iregister_file.vhd:137:9  */
  assign n33806_o = 32'b00000000000000000000000000000111 == n33804_o;
  assign n33807_o = {wr_en1_in, wr_en1_in};
  /* ../../HW/src/ialu/iregister_file.vhd:137:5  */
  assign n33809_o = n33806_o ? n33807_o : 2'b00;
  /* ../../HW/src/ialu/iregister_file.vhd:144:88  */
  assign n33810_o = ~wr_data1_in;
  assign n33811_o = {wr_lane_in, wr_lane_in};
  /* ../../HW/src/ialu/iregister_file.vhd:168:19  */
  assign iregister_ram_i_n33814 = iregister_ram_i_q1_out; // (signal)
  /* ../../HW/src/ialu/iregister_file.vhd:152:1  */
  iregister_ram_5_144 iregister_ram_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .data1_in(wrdata1),
    .rdaddress1_in(rdaddr1),
    .wraddress1_in(wraddr1),
    .wrbyteena1_in(byteena1),
    .wren1_in(n33813_o),
    .rden1_in(rd_en1_in),
    .q1_out(iregister_ram_i_q1_out));
  assign n33826_o = {3'bZ, n33810_o, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in, 3'bZ, wr_data1_in};
  assign n33827_o = {n33811_o, n33809_o, n33802_o, n33795_o, n33788_o, n33781_o, n33774_o, n33767_o, n33760_o};
  /* ../../HW/src/ialu/iregister_file.vhd:122:5  */
  always @(posedge clock_in or posedge n33744_o)
    if (n33744_o)
      n33828_q <= 13'b0000000000000;
    else
      n33828_q <= n33747_o;
  /* ../../HW/src/ialu/iregister_file.vhd:119:1  */
  assign n33829_o = {n33740_o, n33739_o, n33738_o, n33737_o, n33736_o, n33735_o, n33734_o, n33733_o};
endmodule

module xregister_file
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  write_result_vector_in,
   input  [7:0] write_result_lane_in,
   input  [7:0] write_addr_in,
   input  write_result_ena_in,
   input  write_xreg_ena_in,
   input  write_xreg_result_ena_in,
   input  [255:0] write_data_in,
   input  [7:0] write_result_in,
   input  [7:0] read_addr_in,
   output [12:0] read_result_out,
   output [255:0] read_xreg_out);
  wire write_ena;
  wire [271:0] wrdata;
  wire [271:0] q;
  wire [7:0] wraddr;
  wire [7:0] rdaddr;
  wire [33:0] byteena;
  wire [12:0] iregister;
  wire [255:0] read_xreg_r;
  wire [3:0] n33658_o;
  wire [3:0] n33659_o;
  wire [3:0] n33660_o;
  wire [3:0] n33661_o;
  wire [3:0] n33662_o;
  wire [3:0] n33663_o;
  wire [3:0] n33664_o;
  wire [3:0] n33665_o;
  wire [15:0] n33666_o;
  wire [15:0] n33667_o;
  wire [31:0] n33668_o;
  wire [1:0] n33669_o;
  wire [12:0] n33670_o;
  wire n33673_o;
  wire [255:0] n33675_o;
  wire n33682_o;
  wire n33683_o;
  wire n33684_o;
  wire n33685_o;
  wire n33686_o;
  wire n33687_o;
  wire [1:0] n33688_o;
  wire n33689_o;
  wire n33690_o;
  wire n33691_o;
  wire [2:0] n33692_o;
  wire n33693_o;
  wire n33694_o;
  wire n33695_o;
  wire [3:0] n33696_o;
  wire n33697_o;
  wire n33698_o;
  wire n33699_o;
  wire [4:0] n33700_o;
  wire n33701_o;
  wire n33702_o;
  wire n33703_o;
  wire [5:0] n33704_o;
  wire n33705_o;
  wire n33706_o;
  wire n33707_o;
  wire [6:0] n33708_o;
  wire n33709_o;
  wire n33710_o;
  wire n33711_o;
  wire [7:0] n33712_o;
  wire [11:0] n33714_o;
  wire n33715_o;
  wire [12:0] n33716_o;
  wire [12:0] n33717_o;
  wire [12:0] n33718_o;
  wire [271:0] gen2_altsyncram_i_n33720;
  wire [271:0] gen2_altsyncram_i_q_b;
  wire [271:0] n33724_o;
  wire [33:0] n33725_o;
  reg [255:0] n33726_q;
  assign read_result_out = n33670_o;
  assign read_xreg_out = read_xreg_r;
  /* ../../HW/src/pcore/xregister_file.vhd:66:8  */
  assign write_ena = write_xreg_result_ena_in; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:67:8  */
  assign wrdata = n33724_o; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:68:8  */
  assign q = gen2_altsyncram_i_n33720; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:69:8  */
  assign wraddr = write_addr_in; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:70:8  */
  assign rdaddr = read_addr_in; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:71:8  */
  assign byteena = n33725_o; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:72:8  */
  assign iregister = n33718_o; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:73:8  */
  assign read_xreg_r = n33726_q; // (signal)
  /* ../../HW/src/util/arbiter.vhd:74:5  */
  assign n33658_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33659_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33660_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33661_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33662_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33663_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33664_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33665_o = {write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in, write_xreg_ena_in};
  assign n33666_o = {n33658_o, n33659_o, n33660_o, n33661_o};
  assign n33667_o = {n33662_o, n33663_o, n33664_o, n33665_o};
  assign n33668_o = {n33666_o, n33667_o};
  assign n33669_o = {write_result_ena_in, write_result_ena_in};
  /* ../../HW/src/pcore/xregister_file.vhd:85:30  */
  assign n33670_o = q[268:256];
  /* ../../HW/src/pcore/xregister_file.vhd:95:17  */
  assign n33673_o = ~reset_in;
  /* ../../HW/src/pcore/xregister_file.vhd:99:27  */
  assign n33675_o = q[255:0];
  /* ../../HW/src/pcore/xregister_file.vhd:108:46  */
  assign n33682_o = write_result_in[7];
  /* ../../HW/src/pcore/xregister_file.vhd:108:74  */
  assign n33683_o = write_result_lane_in[7];
  /* ../../HW/src/pcore/xregister_file.vhd:108:50  */
  assign n33684_o = n33682_o & n33683_o;
  /* ../../HW/src/pcore/xregister_file.vhd:109:46  */
  assign n33685_o = write_result_in[6];
  /* ../../HW/src/pcore/xregister_file.vhd:109:74  */
  assign n33686_o = write_result_lane_in[6];
  /* ../../HW/src/pcore/xregister_file.vhd:109:50  */
  assign n33687_o = n33685_o & n33686_o;
  /* ../../HW/src/pcore/xregister_file.vhd:108:79  */
  assign n33688_o = {n33684_o, n33687_o};
  /* ../../HW/src/pcore/xregister_file.vhd:110:46  */
  assign n33689_o = write_result_in[5];
  /* ../../HW/src/pcore/xregister_file.vhd:110:74  */
  assign n33690_o = write_result_lane_in[5];
  /* ../../HW/src/pcore/xregister_file.vhd:110:50  */
  assign n33691_o = n33689_o & n33690_o;
  /* ../../HW/src/pcore/xregister_file.vhd:109:79  */
  assign n33692_o = {n33688_o, n33691_o};
  /* ../../HW/src/pcore/xregister_file.vhd:111:46  */
  assign n33693_o = write_result_in[4];
  /* ../../HW/src/pcore/xregister_file.vhd:111:74  */
  assign n33694_o = write_result_lane_in[4];
  /* ../../HW/src/pcore/xregister_file.vhd:111:50  */
  assign n33695_o = n33693_o & n33694_o;
  /* ../../HW/src/pcore/xregister_file.vhd:110:79  */
  assign n33696_o = {n33692_o, n33695_o};
  /* ../../HW/src/pcore/xregister_file.vhd:112:46  */
  assign n33697_o = write_result_in[3];
  /* ../../HW/src/pcore/xregister_file.vhd:112:74  */
  assign n33698_o = write_result_lane_in[3];
  /* ../../HW/src/pcore/xregister_file.vhd:112:50  */
  assign n33699_o = n33697_o & n33698_o;
  /* ../../HW/src/pcore/xregister_file.vhd:111:79  */
  assign n33700_o = {n33696_o, n33699_o};
  /* ../../HW/src/pcore/xregister_file.vhd:113:46  */
  assign n33701_o = write_result_in[2];
  /* ../../HW/src/pcore/xregister_file.vhd:113:74  */
  assign n33702_o = write_result_lane_in[2];
  /* ../../HW/src/pcore/xregister_file.vhd:113:50  */
  assign n33703_o = n33701_o & n33702_o;
  /* ../../HW/src/pcore/xregister_file.vhd:112:79  */
  assign n33704_o = {n33700_o, n33703_o};
  /* ../../HW/src/pcore/xregister_file.vhd:114:46  */
  assign n33705_o = write_result_in[1];
  /* ../../HW/src/pcore/xregister_file.vhd:114:74  */
  assign n33706_o = write_result_lane_in[1];
  /* ../../HW/src/pcore/xregister_file.vhd:114:50  */
  assign n33707_o = n33705_o & n33706_o;
  /* ../../HW/src/pcore/xregister_file.vhd:113:79  */
  assign n33708_o = {n33704_o, n33707_o};
  /* ../../HW/src/pcore/xregister_file.vhd:115:46  */
  assign n33709_o = write_result_in[0];
  /* ../../HW/src/pcore/xregister_file.vhd:115:74  */
  assign n33710_o = write_result_lane_in[0];
  /* ../../HW/src/pcore/xregister_file.vhd:115:50  */
  assign n33711_o = n33709_o & n33710_o;
  /* ../../HW/src/pcore/xregister_file.vhd:114:79  */
  assign n33712_o = {n33708_o, n33711_o};
  /* ../../HW/src/pcore/xregister_file.vhd:118:68  */
  assign n33714_o = write_data_in[12:1];
  /* ../../HW/src/pcore/xregister_file.vhd:119:35  */
  assign n33715_o = write_result_in[0];
  assign n33716_o = {n33714_o, n33715_o};
  assign n33717_o = {5'b00000, n33712_o};
  /* ../../HW/src/pcore/xregister_file.vhd:107:1  */
  assign n33718_o = write_result_vector_in ? n33717_o : n33716_o;
  /* ../../HW/src/pcore/xregister_file.vhd:164:16  */
  assign gen2_altsyncram_i_n33720 = gen2_altsyncram_i_q_b; // (signal)
  /* ../../HW/src/pcore/xregister_file.vhd:147:1  */
  ramw_256_256_8_8_272_272 gen2_altsyncram_i (
    .clock(clock_in),
    .clock_x2(clock_x2_in),
    .address_a(wraddr),
    .byteena_a(byteena),
    .data_a(wrdata),
    .wren_a(write_ena),
    .address_b(rdaddr),
    .q_b(gen2_altsyncram_i_q_b));
  assign n33724_o = {3'bZ, iregister, write_data_in};
  assign n33725_o = {n33669_o, n33668_o};
  /* ../../HW/src/pcore/xregister_file.vhd:98:8  */
  always @(posedge clock_in or posedge n33673_o)
    if (n33673_o)
      n33726_q <= 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n33726_q <= n33675_o;
endmodule

module arbiter_16_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clock_in,
   input  reset_in,
   input  [15:0] req_in,
   output [15:0] gnt_out,
   output gnt_valid_out);
  wire [15:0] gnt_r;
  wire [15:0] gnt;
  wire [15:0] gnt1;
  wire [15:0] gnt2;
  wire [15:0] req;
  wire [15:0] n33619_o;
  wire [15:0] n33620_o;
  wire [15:0] n33621_o;
  wire [15:0] n33622_o;
  wire [15:0] n33623_o;
  wire n33625_o;
  wire [15:0] n33626_o;
  wire n33629_o;
  wire n33630_o;
  wire n33635_o;
  wire n33638_o;
  wire [15:0] n33640_o;
  wire [15:0] n33641_o;
  wire [15:0] n33642_o;
  wire [15:0] n33654_o;
  reg [15:0] n33655_q;
  assign gnt_out = gnt2;
  assign gnt_valid_out = n33630_o;
  /* ../../HW/src/util/arbiter.vhd:45:8  */
  assign gnt_r = n33655_q; // (signal)
  /* ../../HW/src/util/arbiter.vhd:46:8  */
  assign gnt = n33620_o; // (signal)
  /* ../../HW/src/util/arbiter.vhd:47:8  */
  assign gnt1 = n33623_o; // (signal)
  /* ../../HW/src/util/arbiter.vhd:48:8  */
  assign gnt2 = n33626_o; // (signal)
  /* ../../HW/src/util/arbiter.vhd:49:8  */
  assign req = n33621_o; // (signal)
  /* ../../HW/src/util/arbiter.vhd:60:36  */
  assign n33619_o = -req_in;
  /* ../../HW/src/util/arbiter.vhd:60:15  */
  assign n33620_o = req_in & n33619_o;
  /* ../../HW/src/util/arbiter.vhd:61:15  */
  assign n33621_o = req_in & gnt_r;
  /* ../../HW/src/util/arbiter.vhd:62:34  */
  assign n33622_o = -req;
  /* ../../HW/src/util/arbiter.vhd:62:13  */
  assign n33623_o = req & n33622_o;
  /* ../../HW/src/util/arbiter.vhd:63:23  */
  assign n33625_o = req != 16'b0000000000000000;
  /* ../../HW/src/util/arbiter.vhd:63:14  */
  assign n33626_o = n33625_o ? gnt1 : gnt;
  /* ../../HW/src/util/arbiter.vhd:65:33  */
  assign n33629_o = req_in == 16'b0000000000000000;
  /* ../../HW/src/util/arbiter.vhd:65:22  */
  assign n33630_o = n33629_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/arbiter.vhd:74:17  */
  assign n33635_o = ~reset_in;
  /* ../../HW/src/util/arbiter.vhd:79:23  */
  assign n33638_o = req_in != 16'b0000000000000000;
  /* ../../HW/src/util/arbiter.vhd:80:64  */
  assign n33640_o = gnt2 - 16'b0000000000000001;
  /* ../../HW/src/util/arbiter.vhd:80:69  */
  assign n33641_o = n33640_o | gnt2;
  /* ../../HW/src/util/arbiter.vhd:80:27  */
  assign n33642_o = ~n33641_o;
  /* ../../HW/src/util/arbiter.vhd:77:9  */
  assign n33654_o = n33638_o ? n33642_o : gnt_r;
  /* ../../HW/src/util/arbiter.vhd:77:9  */
  always @(posedge clock_in or posedge n33635_o)
    if (n33635_o)
      n33655_q <= 16'b0000000000000000;
    else
      n33655_q <= n33654_o;
endmodule

module delayv_16_1
  (input  clock_in,
   input  reset_in,
   input  [15:0] in_in,
   input  enable_in,
   output [15:0] out_out);
  wire [15:0] fifo_r;
  wire n33608_o;
  wire [15:0] n33615_o;
  reg [15:0] n33616_q;
  assign out_out = fifo_r;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n33616_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n33608_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:56:9  */
  assign n33615_o = enable_in ? in_in : fifo_r;
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n33608_o)
    if (n33608_o)
      n33616_q <= 16'b0000000000000000;
    else
      n33616_q <= n33615_o;
endmodule

module spram_be_1024_10_128
  (input  [9:0] address_a,
   input  clock0,
   input  [127:0] data_a,
   input  wren_a,
   input  [15:0] byteena_a,
   output [127:0] q_a);
  wire [127:0] q;
  wire [127:0] data;
  wire [9:0] address_r;
  wire [7:0] n33369_o;
  wire [7:0] n33370_o;
  wire [7:0] n33371_o;
  wire [7:0] n33372_o;
  wire [7:0] n33373_o;
  wire [7:0] n33374_o;
  wire [7:0] n33375_o;
  wire [7:0] n33376_o;
  wire [7:0] n33377_o;
  wire [7:0] n33378_o;
  wire [7:0] n33379_o;
  wire [7:0] n33380_o;
  wire [7:0] n33381_o;
  wire [7:0] n33382_o;
  wire [7:0] n33383_o;
  wire [7:0] n33384_o;
  wire [7:0] n33385_o;
  wire [7:0] n33386_o;
  wire [7:0] n33387_o;
  wire [7:0] n33388_o;
  wire [7:0] n33389_o;
  wire [7:0] n33390_o;
  wire [7:0] n33391_o;
  wire [7:0] n33392_o;
  wire [7:0] n33393_o;
  wire [7:0] n33394_o;
  wire [7:0] n33395_o;
  wire [7:0] n33396_o;
  wire [7:0] n33397_o;
  wire [7:0] n33398_o;
  wire [7:0] n33399_o;
  wire [7:0] n33400_o;
  wire n33404_o;
  wire [7:0] n33409_o;
  wire n33412_o;
  wire [7:0] n33417_o;
  wire n33420_o;
  wire [7:0] n33425_o;
  wire n33428_o;
  wire [7:0] n33433_o;
  wire n33436_o;
  wire [7:0] n33441_o;
  wire n33444_o;
  wire [7:0] n33449_o;
  wire n33452_o;
  wire [7:0] n33457_o;
  wire n33460_o;
  wire [7:0] n33465_o;
  wire n33468_o;
  wire [7:0] n33473_o;
  wire n33476_o;
  wire [7:0] n33481_o;
  wire n33484_o;
  wire [7:0] n33489_o;
  wire n33492_o;
  wire [7:0] n33497_o;
  wire n33500_o;
  wire [7:0] n33505_o;
  wire n33508_o;
  wire [7:0] n33513_o;
  wire n33516_o;
  wire [7:0] n33521_o;
  wire n33524_o;
  wire [7:0] n33529_o;
  wire n33536_o;
  wire n33538_o;
  wire n33540_o;
  wire n33542_o;
  wire n33544_o;
  wire n33546_o;
  wire n33548_o;
  wire n33550_o;
  wire n33552_o;
  wire n33554_o;
  wire n33556_o;
  wire n33558_o;
  wire n33560_o;
  wire n33562_o;
  wire n33564_o;
  wire n33566_o;
  wire [127:0] n33569_o;
  reg [9:0] n33570_q;
  wire [127:0] n33571_o;
  wire [7:0] n33572_data; // mem_rd
  wire [7:0] n33573_data; // mem_rd
  wire [7:0] n33574_data; // mem_rd
  wire [7:0] n33575_data; // mem_rd
  wire [7:0] n33576_data; // mem_rd
  wire [7:0] n33577_data; // mem_rd
  wire [7:0] n33578_data; // mem_rd
  wire [7:0] n33579_data; // mem_rd
  wire [7:0] n33580_data; // mem_rd
  wire [7:0] n33581_data; // mem_rd
  wire [7:0] n33582_data; // mem_rd
  wire [7:0] n33583_data; // mem_rd
  wire [7:0] n33584_data; // mem_rd
  wire [7:0] n33585_data; // mem_rd
  wire [7:0] n33586_data; // mem_rd
  wire [7:0] n33587_data; // mem_rd
  wire [127:0] n33588_o;
  assign q_a = n33571_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:51:8  */
  assign q = n33588_o; // (signal)
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:52:8  */
  assign data = n33569_o; // (signal)
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:53:8  */
  assign address_r = n33570_q; // (signal)
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33369_o = q[127:120];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33370_o = q[119:112];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33371_o = q[111:104];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33372_o = q[103:96];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33373_o = q[95:88];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33374_o = q[87:80];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33375_o = q[79:72];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33376_o = q[71:64];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33377_o = q[63:56];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33378_o = q[55:48];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33379_o = q[47:40];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33380_o = q[39:32];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33381_o = q[31:24];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33382_o = q[23:16];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33383_o = q[15:8];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:61:30  */
  assign n33384_o = q[7:0];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33385_o = data_a[7:0];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33386_o = data_a[15:8];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33387_o = data_a[23:16];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33388_o = data_a[31:24];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33389_o = data_a[39:32];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33390_o = data_a[47:40];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33391_o = data_a[55:48];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33392_o = data_a[63:56];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33393_o = data_a[71:64];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33394_o = data_a[79:72];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33395_o = data_a[87:80];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33396_o = data_a[95:88];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33397_o = data_a[103:96];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33398_o = data_a[111:104];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33399_o = data_a[119:112];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:65:21  */
  assign n33400_o = data_a[127:120];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33404_o = byteena_a[0];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33409_o = data[127:120];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33412_o = byteena_a[1];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33417_o = data[119:112];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33420_o = byteena_a[2];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33425_o = data[111:104];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33428_o = byteena_a[3];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33433_o = data[103:96];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33436_o = byteena_a[4];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33441_o = data[95:88];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33444_o = byteena_a[5];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33449_o = data[87:80];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33452_o = byteena_a[6];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33457_o = data[79:72];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33460_o = byteena_a[7];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33465_o = data[71:64];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33468_o = byteena_a[8];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33473_o = data[63:56];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33476_o = byteena_a[9];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33481_o = data[55:48];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33484_o = byteena_a[10];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33489_o = data[47:40];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33492_o = byteena_a[11];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33497_o = data[39:32];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33500_o = byteena_a[12];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33505_o = data[31:24];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33508_o = byteena_a[13];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33513_o = data[23:16];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33516_o = byteena_a[14];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33521_o = data[15:8];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:73:25  */
  assign n33524_o = byteena_a[15];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:69  */
  assign n33529_o = data[7:0];
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33536_o = wren_a & n33524_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33538_o = wren_a & n33516_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33540_o = wren_a & n33508_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33542_o = wren_a & n33500_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33544_o = wren_a & n33492_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33546_o = wren_a & n33484_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33548_o = wren_a & n33476_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33550_o = wren_a & n33468_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33552_o = wren_a & n33460_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33554_o = wren_a & n33452_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33556_o = wren_a & n33444_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33558_o = wren_a & n33436_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33560_o = wren_a & n33428_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33562_o = wren_a & n33420_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33564_o = wren_a & n33412_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:30:8  */
  assign n33566_o = wren_a & n33404_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:70:4  */
  assign n33569_o = {n33385_o, n33386_o, n33387_o, n33388_o, n33389_o, n33390_o, n33391_o, n33392_o, n33393_o, n33394_o, n33395_o, n33396_o, n33397_o, n33398_o, n33399_o, n33400_o};
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:70:4  */
  always @(posedge clock0)
    n33570_q <= address_a;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:70:4  */
  assign n33571_o = {n33384_o, n33383_o, n33382_o, n33381_o, n33380_o, n33379_o, n33378_o, n33377_o, n33376_o, n33375_o, n33374_o, n33373_o, n33372_o, n33371_o, n33370_o, n33369_o};
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:59:16  */
  reg [7:0] ram_block_n1[1023:0] ; // memory
  assign n33572_data = ram_block_n1[address_r];
  always @(posedge clock0)
    if (n33536_o)
      ram_block_n1[address_a] <= n33529_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:59:16  */
  reg [7:0] ram_block_n2[1023:0] ; // memory
  assign n33573_data = ram_block_n2[address_r];
  always @(posedge clock0)
    if (n33538_o)
      ram_block_n2[address_a] <= n33521_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n3[1023:0] ; // memory
  assign n33574_data = ram_block_n3[address_r];
  always @(posedge clock0)
    if (n33540_o)
      ram_block_n3[address_a] <= n33513_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n4[1023:0] ; // memory
  assign n33575_data = ram_block_n4[address_r];
  always @(posedge clock0)
    if (n33542_o)
      ram_block_n4[address_a] <= n33505_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n5[1023:0] ; // memory
  assign n33576_data = ram_block_n5[address_r];
  always @(posedge clock0)
    if (n33544_o)
      ram_block_n5[address_a] <= n33497_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n6[1023:0] ; // memory
  assign n33577_data = ram_block_n6[address_r];
  always @(posedge clock0)
    if (n33546_o)
      ram_block_n6[address_a] <= n33489_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n7[1023:0] ; // memory
  assign n33578_data = ram_block_n7[address_r];
  always @(posedge clock0)
    if (n33548_o)
      ram_block_n7[address_a] <= n33481_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n8[1023:0] ; // memory
  assign n33579_data = ram_block_n8[address_r];
  always @(posedge clock0)
    if (n33550_o)
      ram_block_n8[address_a] <= n33473_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n9[1023:0] ; // memory
  assign n33580_data = ram_block_n9[address_r];
  always @(posedge clock0)
    if (n33552_o)
      ram_block_n9[address_a] <= n33465_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n10[1023:0] ; // memory
  assign n33581_data = ram_block_n10[address_r];
  always @(posedge clock0)
    if (n33554_o)
      ram_block_n10[address_a] <= n33457_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n11[1023:0] ; // memory
  assign n33582_data = ram_block_n11[address_r];
  always @(posedge clock0)
    if (n33556_o)
      ram_block_n11[address_a] <= n33449_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n12[1023:0] ; // memory
  assign n33583_data = ram_block_n12[address_r];
  always @(posedge clock0)
    if (n33558_o)
      ram_block_n12[address_a] <= n33441_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n13[1023:0] ; // memory
  assign n33584_data = ram_block_n13[address_r];
  always @(posedge clock0)
    if (n33560_o)
      ram_block_n13[address_a] <= n33433_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n14[1023:0] ; // memory
  assign n33585_data = ram_block_n14[address_r];
  always @(posedge clock0)
    if (n33562_o)
      ram_block_n14[address_a] <= n33425_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n15[1023:0] ; // memory
  assign n33586_data = ram_block_n15[address_r];
  always @(posedge clock0)
    if (n33564_o)
      ram_block_n15[address_a] <= n33417_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  reg [7:0] ram_block_n16[1023:0] ; // memory
  assign n33587_data = ram_block_n16[address_r];
  always @(posedge clock0)
    if (n33566_o)
      ram_block_n16[address_a] <= n33409_o;
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:59:16  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  assign n33588_o = {n33587_data, n33586_data, n33585_data, n33584_data, n33583_data, n33582_data, n33581_data, n33580_data, n33579_data, n33578_data, n33577_data, n33576_data, n33575_data, n33574_data, n33573_data, n33572_data};
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
  /* ../../HW/platform/simulation/SPRAM_BE.vhd:74:26  */
endmodule

module scfifo_64_9_1_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clock_in,
   input  reset_in,
   input  [63:0] data_in,
   input  write_in,
   input  read_in,
   output [63:0] q_out,
   output [8:0] ravail_out,
   output [8:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [63:0] q;
  wire [63:0] q_r;
  wire [8:0] address_a;
  wire [8:0] address_b;
  wire [8:0] waddr_r;
  wire [8:0] waddr_rr;
  wire [8:0] raddr_r;
  wire [8:0] raddr;
  wire [8:0] ravail;
  wire [8:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [63:0] ram_i_n33296;
  wire [63:0] ram_i_q_b;
  wire [8:0] n33299_o;
  wire [8:0] n33300_o;
  wire n33301_o;
  wire n33304_o;
  wire n33305_o;
  wire [8:0] n33308_o;
  wire [8:0] n33309_o;
  wire n33312_o;
  wire [8:0] n33315_o;
  wire [8:0] n33317_o;
  wire n33318_o;
  wire n33321_o;
  wire [8:0] n33323_o;
  wire n33324_o;
  wire n33327_o;
  wire n33329_o;
  wire n33331_o;
  wire n33334_o;
  wire [63:0] n33354_o;
  reg [63:0] n33355_q;
  wire [8:0] n33356_o;
  reg [8:0] n33357_q;
  reg [8:0] n33358_q;
  reg [8:0] n33359_q;
  reg n33361_q;
  reg n33362_q;
  assign q_out = q_r;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n33301_o;
  assign full_out = full_r;
  assign almost_full_out = n33305_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n33296; // (signal)
  /* ../../HW/src/util/fifo.vhd:54:8  */
  assign q_r = n33355_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n33357_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n33358_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n33359_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n33309_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n33299_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n33300_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n33361_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n33362_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n33296 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_512_512_9_9_64_64 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n33299_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n33300_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n33301_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n33304_o = $unsigned(wused) >= $unsigned(9'b000000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n33305_o = n33304_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n33308_o = raddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n33309_o = read_in ? n33308_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n33312_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n33315_o = waddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n33317_o = waddr_r + 9'b000000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n33318_o = n33317_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n33321_o = n33318_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n33323_o = waddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n33324_o = n33323_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n33327_o = n33324_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n33329_o = write_in ? n33321_o : n33327_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n33331_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n33334_o = n33331_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n33354_o = read_in ? q : q_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33312_o)
    if (n33312_o)
      n33355_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n33355_q <= n33354_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n33356_o = write_in ? n33315_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33312_o)
    if (n33312_o)
      n33357_q <= 9'b000000000;
    else
      n33357_q <= n33356_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33312_o)
    if (n33312_o)
      n33358_q <= 9'b000000000;
    else
      n33358_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33312_o)
    if (n33312_o)
      n33359_q <= 9'b000000000;
    else
      n33359_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33312_o)
    if (n33312_o)
      n33361_q <= 1'b0;
    else
      n33361_q <= n33334_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33312_o)
    if (n33312_o)
      n33362_q <= 1'b0;
    else
      n33362_q <= n33329_o;
endmodule

module scfifo_132_9_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [131:0] data_in,
   input  write_in,
   input  read_in,
   output [131:0] q_out,
   output [8:0] ravail_out,
   output [8:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [131:0] q;
  wire [8:0] address_a;
  wire [8:0] address_b;
  wire [8:0] waddr_r;
  wire [8:0] waddr_rr;
  wire [8:0] raddr_r;
  wire [8:0] raddr;
  wire [8:0] ravail;
  wire [8:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [131:0] ram_i_n33223;
  wire [131:0] ram_i_q_b;
  wire [8:0] n33226_o;
  wire [8:0] n33227_o;
  wire n33228_o;
  wire n33231_o;
  wire n33232_o;
  wire [8:0] n33235_o;
  wire [8:0] n33236_o;
  wire n33239_o;
  wire [8:0] n33242_o;
  wire [8:0] n33244_o;
  wire n33245_o;
  wire n33248_o;
  wire [8:0] n33250_o;
  wire n33251_o;
  wire n33254_o;
  wire n33256_o;
  wire n33258_o;
  wire n33261_o;
  wire [8:0] n33283_o;
  reg [8:0] n33284_q;
  reg [8:0] n33285_q;
  reg [8:0] n33286_q;
  reg n33288_q;
  reg n33289_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n33228_o;
  assign full_out = full_r;
  assign almost_full_out = n33232_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n33223; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n33284_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n33285_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n33286_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n33236_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n33226_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n33227_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n33288_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n33289_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n33223 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_512_512_9_9_132_132 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n33226_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n33227_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n33228_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n33231_o = $unsigned(wused) >= $unsigned(9'b000000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n33232_o = n33231_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n33235_o = raddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n33236_o = read_in ? n33235_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n33239_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n33242_o = waddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n33244_o = waddr_r + 9'b000000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n33245_o = n33244_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n33248_o = n33245_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n33250_o = waddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n33251_o = n33250_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n33254_o = n33251_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n33256_o = write_in ? n33248_o : n33254_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n33258_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n33261_o = n33258_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n33283_o = write_in ? n33242_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33239_o)
    if (n33239_o)
      n33284_q <= 9'b000000000;
    else
      n33284_q <= n33283_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33239_o)
    if (n33239_o)
      n33285_q <= 9'b000000000;
    else
      n33285_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33239_o)
    if (n33239_o)
      n33286_q <= 9'b000000000;
    else
      n33286_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33239_o)
    if (n33239_o)
      n33288_q <= 1'b0;
    else
      n33288_q <= n33261_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n33239_o)
    if (n33239_o)
      n33289_q <= 1'b0;
    else
      n33289_q <= n33256_o;
endmodule

module delayv_64_7
  (input  clock_in,
   input  reset_in,
   input  [63:0] in_in,
   input  enable_in,
   output [63:0] out_out);
  wire [447:0] fifo_r;
  wire [63:0] n33179_o;
  wire n33182_o;
  wire [63:0] n33191_o;
  wire [63:0] n33192_o;
  wire [63:0] n33193_o;
  wire [63:0] n33194_o;
  wire [63:0] n33195_o;
  wire [63:0] n33196_o;
  wire [63:0] n33197_o;
  wire [63:0] n33198_o;
  wire [63:0] n33199_o;
  wire [63:0] n33200_o;
  wire [63:0] n33201_o;
  wire [63:0] n33202_o;
  wire [63:0] n33203_o;
  wire [63:0] n33204_o;
  wire [63:0] n33205_o;
  wire [63:0] n33206_o;
  wire [63:0] n33207_o;
  wire [63:0] n33208_o;
  wire [63:0] n33209_o;
  wire [63:0] n33210_o;
  wire [447:0] n33211_o;
  wire [447:0] n33213_o;
  reg [447:0] n33216_q;
  assign out_out = n33179_o;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n33216_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:48:18  */
  assign n33179_o = fifo_r[63:0];
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n33182_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33191_o = fifo_r[127:64];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33192_o = fifo_r[63:0];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33193_o = enable_in ? n33191_o : n33192_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33194_o = fifo_r[191:128];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33195_o = fifo_r[127:64];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33196_o = enable_in ? n33194_o : n33195_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33197_o = fifo_r[255:192];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33198_o = fifo_r[191:128];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33199_o = enable_in ? n33197_o : n33198_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33200_o = fifo_r[319:256];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33201_o = fifo_r[255:192];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33202_o = enable_in ? n33200_o : n33201_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33203_o = fifo_r[383:320];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33204_o = fifo_r[319:256];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33205_o = enable_in ? n33203_o : n33204_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33206_o = fifo_r[447:384];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33207_o = fifo_r[383:320];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33208_o = enable_in ? n33206_o : n33207_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33209_o = fifo_r[447:384];
  /* ../../HW/src/util/delayv.vhd:64:13  */
  assign n33210_o = enable_in ? in_in : n33209_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33211_o = {n33210_o, n33208_o, n33205_o, n33202_o, n33199_o, n33196_o, n33193_o};
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33213_o = {64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n33182_o)
    if (n33182_o)
      n33216_q <= n33213_o;
    else
      n33216_q <= n33211_o;
endmodule

module delayv_64_4
  (input  clock_in,
   input  reset_in,
   input  [63:0] in_in,
   input  enable_in,
   output [63:0] out_out);
  wire [255:0] fifo_r;
  wire [63:0] n33152_o;
  wire n33155_o;
  wire [63:0] n33161_o;
  wire [63:0] n33162_o;
  wire [63:0] n33163_o;
  wire [63:0] n33164_o;
  wire [63:0] n33165_o;
  wire [63:0] n33166_o;
  wire [63:0] n33167_o;
  wire [63:0] n33168_o;
  wire [63:0] n33169_o;
  wire [63:0] n33170_o;
  wire [63:0] n33171_o;
  wire [255:0] n33172_o;
  wire [255:0] n33174_o;
  reg [255:0] n33177_q;
  assign out_out = n33152_o;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n33177_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:48:18  */
  assign n33152_o = fifo_r[63:0];
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n33155_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33161_o = fifo_r[127:64];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33162_o = fifo_r[63:0];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33163_o = enable_in ? n33161_o : n33162_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33164_o = fifo_r[191:128];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33165_o = fifo_r[127:64];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33166_o = enable_in ? n33164_o : n33165_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33167_o = fifo_r[255:192];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33168_o = fifo_r[191:128];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33169_o = enable_in ? n33167_o : n33168_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33170_o = fifo_r[255:192];
  /* ../../HW/src/util/delayv.vhd:64:13  */
  assign n33171_o = enable_in ? in_in : n33170_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33172_o = {n33171_o, n33169_o, n33166_o, n33163_o};
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33174_o = {64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n33155_o)
    if (n33155_o)
      n33177_q <= n33174_o;
    else
      n33177_q <= n33172_o;
endmodule

module delayv_64_8
  (input  clock_in,
   input  reset_in,
   input  [63:0] in_in,
   input  enable_in,
   output [63:0] out_out);
  wire [511:0] fifo_r;
  wire [63:0] n33109_o;
  wire n33112_o;
  wire [63:0] n33122_o;
  wire [63:0] n33123_o;
  wire [63:0] n33124_o;
  wire [63:0] n33125_o;
  wire [63:0] n33126_o;
  wire [63:0] n33127_o;
  wire [63:0] n33128_o;
  wire [63:0] n33129_o;
  wire [63:0] n33130_o;
  wire [63:0] n33131_o;
  wire [63:0] n33132_o;
  wire [63:0] n33133_o;
  wire [63:0] n33134_o;
  wire [63:0] n33135_o;
  wire [63:0] n33136_o;
  wire [63:0] n33137_o;
  wire [63:0] n33138_o;
  wire [63:0] n33139_o;
  wire [63:0] n33140_o;
  wire [63:0] n33141_o;
  wire [63:0] n33142_o;
  wire [63:0] n33143_o;
  wire [63:0] n33144_o;
  wire [511:0] n33145_o;
  wire [511:0] n33147_o;
  reg [511:0] n33150_q;
  assign out_out = n33109_o;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n33150_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:48:18  */
  assign n33109_o = fifo_r[63:0];
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n33112_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33122_o = fifo_r[127:64];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33123_o = fifo_r[63:0];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33124_o = enable_in ? n33122_o : n33123_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33125_o = fifo_r[191:128];
  /* ../../HW/src/dp/dp_gen.vhd:766:1  */
  assign n33126_o = fifo_r[127:64];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33127_o = enable_in ? n33125_o : n33126_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33128_o = fifo_r[255:192];
  /* ../../HW/src/dp/dp_gen.vhd:766:1  */
  assign n33129_o = fifo_r[191:128];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33130_o = enable_in ? n33128_o : n33129_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33131_o = fifo_r[319:256];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33132_o = fifo_r[255:192];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33133_o = enable_in ? n33131_o : n33132_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33134_o = fifo_r[383:320];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33135_o = fifo_r[319:256];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33136_o = enable_in ? n33134_o : n33135_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33137_o = fifo_r[447:384];
  /* ../../HW/src/dp/dp_gen.vhd:766:1  */
  assign n33138_o = fifo_r[383:320];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33139_o = enable_in ? n33137_o : n33138_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33140_o = fifo_r[511:448];
  assign n33141_o = fifo_r[447:384];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33142_o = enable_in ? n33140_o : n33141_o;
  assign n33143_o = fifo_r[511:448];
  /* ../../HW/src/util/delayv.vhd:64:13  */
  assign n33144_o = enable_in ? in_in : n33143_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33145_o = {n33144_o, n33142_o, n33139_o, n33136_o, n33133_o, n33130_o, n33127_o, n33124_o};
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33147_o = {64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000, 64'b0000000000000000000000000000000000000000000000000000000000000000};
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n33112_o)
    if (n33112_o)
      n33150_q <= n33147_o;
    else
      n33150_q <= n33145_o;
endmodule

module delayv_6_8
  (input  clock_in,
   input  reset_in,
   input  [5:0] in_in,
   input  enable_in,
   output [5:0] out_out);
  wire [47:0] fifo_r;
  wire [5:0] n33066_o;
  wire n33069_o;
  wire [5:0] n33079_o;
  wire [5:0] n33080_o;
  wire [5:0] n33081_o;
  wire [5:0] n33082_o;
  wire [5:0] n33083_o;
  wire [5:0] n33084_o;
  wire [5:0] n33085_o;
  wire [5:0] n33086_o;
  wire [5:0] n33087_o;
  wire [5:0] n33088_o;
  wire [5:0] n33089_o;
  wire [5:0] n33090_o;
  wire [5:0] n33091_o;
  wire [5:0] n33092_o;
  wire [5:0] n33093_o;
  wire [5:0] n33094_o;
  wire [5:0] n33095_o;
  wire [5:0] n33096_o;
  wire [5:0] n33097_o;
  wire [5:0] n33098_o;
  wire [5:0] n33099_o;
  wire [5:0] n33100_o;
  wire [5:0] n33101_o;
  wire [47:0] n33102_o;
  wire [47:0] n33104_o;
  reg [47:0] n33107_q;
  assign out_out = n33066_o;
  /* ../../HW/src/util/delayv.vhd:46:8  */
  assign fifo_r = n33107_q; // (signal)
  /* ../../HW/src/util/delayv.vhd:48:18  */
  assign n33066_o = fifo_r[5:0];
  /* ../../HW/src/util/delayv.vhd:51:16  */
  assign n33069_o = ~reset_in;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33079_o = fifo_r[11:6];
  /* ../../HW/src/dp/dp_gen.vhd:1800:49  */
  assign n33080_o = fifo_r[5:0];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33081_o = enable_in ? n33079_o : n33080_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33082_o = fifo_r[17:12];
  /* ../../HW/src/dp/dp_gen.vhd:1752:49  */
  assign n33083_o = fifo_r[11:6];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33084_o = enable_in ? n33082_o : n33083_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33085_o = fifo_r[23:18];
  assign n33086_o = fifo_r[17:12];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33087_o = enable_in ? n33085_o : n33086_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33088_o = fifo_r[29:24];
  assign n33089_o = fifo_r[23:18];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33090_o = enable_in ? n33088_o : n33089_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33091_o = fifo_r[35:30];
  assign n33092_o = fifo_r[29:24];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33093_o = enable_in ? n33091_o : n33092_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33094_o = fifo_r[41:36];
  assign n33095_o = fifo_r[35:30];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33096_o = enable_in ? n33094_o : n33095_o;
  /* ../../HW/src/util/delayv.vhd:60:44  */
  assign n33097_o = fifo_r[47:42];
  assign n33098_o = fifo_r[41:36];
  /* ../../HW/src/util/delayv.vhd:59:21  */
  assign n33099_o = enable_in ? n33097_o : n33098_o;
  assign n33100_o = fifo_r[47:42];
  /* ../../HW/src/util/delayv.vhd:64:13  */
  assign n33101_o = enable_in ? in_in : n33100_o;
  /* ../../HW/src/dp/dp_gen.vhd:776:5  */
  assign n33102_o = {n33101_o, n33099_o, n33096_o, n33093_o, n33090_o, n33087_o, n33084_o, n33081_o};
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n33104_o = {6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000};
  /* ../../HW/src/util/delayv.vhd:56:9  */
  always @(posedge clock_in or posedge n33069_o)
    if (n33069_o)
      n33107_q <= n33104_o;
    else
      n33107_q <= n33102_o;
endmodule

module delayi_5_8
  (input  clock_in,
   input  reset_in,
   input  [4:0] in_in,
   input  enable_in,
   output [4:0] out_out);
  wire [39:0] fifo_r;
  wire [4:0] n33023_o;
  wire n33026_o;
  wire [4:0] n33036_o;
  wire [4:0] n33037_o;
  wire [4:0] n33038_o;
  wire [4:0] n33039_o;
  wire [4:0] n33040_o;
  wire [4:0] n33041_o;
  wire [4:0] n33042_o;
  wire [4:0] n33043_o;
  wire [4:0] n33044_o;
  wire [4:0] n33045_o;
  wire [4:0] n33046_o;
  wire [4:0] n33047_o;
  wire [4:0] n33048_o;
  wire [4:0] n33049_o;
  wire [4:0] n33050_o;
  wire [4:0] n33051_o;
  wire [4:0] n33052_o;
  wire [4:0] n33053_o;
  wire [4:0] n33054_o;
  wire [4:0] n33055_o;
  wire [4:0] n33056_o;
  wire [4:0] n33057_o;
  wire [4:0] n33058_o;
  wire [39:0] n33059_o;
  wire [39:0] n33061_o;
  reg [39:0] n33064_q;
  assign out_out = n33023_o;
  /* ../../HW/src/util/delayi.vhd:46:8  */
  assign fifo_r = n33064_q; // (signal)
  /* ../../HW/src/util/delayi.vhd:48:18  */
  assign n33023_o = fifo_r[4:0];
  /* ../../HW/src/util/delayi.vhd:51:16  */
  assign n33026_o = ~reset_in;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33036_o = fifo_r[9:5];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n33037_o = fifo_r[4:0];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33038_o = enable_in ? n33036_o : n33037_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33039_o = fifo_r[14:10];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n33040_o = fifo_r[9:5];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33041_o = enable_in ? n33039_o : n33040_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33042_o = fifo_r[19:15];
  assign n33043_o = fifo_r[14:10];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33044_o = enable_in ? n33042_o : n33043_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33045_o = fifo_r[24:20];
  assign n33046_o = fifo_r[19:15];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33047_o = enable_in ? n33045_o : n33046_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33048_o = fifo_r[29:25];
  assign n33049_o = fifo_r[24:20];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33050_o = enable_in ? n33048_o : n33049_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33051_o = fifo_r[34:30];
  assign n33052_o = fifo_r[29:25];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33053_o = enable_in ? n33051_o : n33052_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33054_o = fifo_r[39:35];
  assign n33055_o = fifo_r[34:30];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33056_o = enable_in ? n33054_o : n33055_o;
  assign n33057_o = fifo_r[39:35];
  /* ../../HW/src/util/delayi.vhd:64:13  */
  assign n33058_o = enable_in ? in_in : n33057_o;
  assign n33059_o = {n33058_o, n33056_o, n33053_o, n33050_o, n33047_o, n33044_o, n33041_o, n33038_o};
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n33061_o = {5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000};
  /* ../../HW/src/util/delayi.vhd:56:9  */
  always @(posedge clock_in or posedge n33026_o)
    if (n33026_o)
      n33064_q <= n33061_o;
    else
      n33064_q <= n33059_o;
endmodule

module delayi_1_8
  (input  clock_in,
   input  reset_in,
   input  in_in,
   input  enable_in,
   output out_out);
  wire [7:0] fifo_r;
  wire n32980_o;
  wire n32983_o;
  wire n32993_o;
  wire n32994_o;
  wire n32995_o;
  wire n32996_o;
  wire n32997_o;
  wire n32998_o;
  wire n32999_o;
  wire n33000_o;
  wire n33001_o;
  wire n33002_o;
  wire n33003_o;
  wire n33004_o;
  wire n33005_o;
  wire n33006_o;
  wire n33007_o;
  wire n33008_o;
  wire n33009_o;
  wire n33010_o;
  wire n33011_o;
  wire n33012_o;
  wire n33013_o;
  wire n33014_o;
  wire n33015_o;
  wire [7:0] n33016_o;
  wire [7:0] n33018_o;
  reg [7:0] n33021_q;
  assign out_out = n32980_o;
  /* ../../HW/src/util/delayi.vhd:46:8  */
  assign fifo_r = n33021_q; // (signal)
  /* ../../HW/src/util/delayi.vhd:48:18  */
  assign n32980_o = fifo_r[0];
  /* ../../HW/src/util/delayi.vhd:51:16  */
  assign n32983_o = ~reset_in;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32993_o = fifo_r[1];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32994_o = fifo_r[0];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32995_o = enable_in ? n32993_o : n32994_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32996_o = fifo_r[2];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32997_o = fifo_r[1];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32998_o = enable_in ? n32996_o : n32997_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32999_o = fifo_r[3];
  assign n33000_o = fifo_r[2];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33001_o = enable_in ? n32999_o : n33000_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33002_o = fifo_r[4];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n33003_o = fifo_r[3];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33004_o = enable_in ? n33002_o : n33003_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33005_o = fifo_r[5];
  assign n33006_o = fifo_r[4];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33007_o = enable_in ? n33005_o : n33006_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33008_o = fifo_r[6];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n33009_o = fifo_r[5];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33010_o = enable_in ? n33008_o : n33009_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n33011_o = fifo_r[7];
  assign n33012_o = fifo_r[6];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n33013_o = enable_in ? n33011_o : n33012_o;
  assign n33014_o = fifo_r[7];
  /* ../../HW/src/util/delayi.vhd:64:13  */
  assign n33015_o = enable_in ? in_in : n33014_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n33016_o = {n33015_o, n33013_o, n33010_o, n33007_o, n33004_o, n33001_o, n32998_o, n32995_o};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n33018_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/util/delayi.vhd:56:9  */
  always @(posedge clock_in or posedge n32983_o)
    if (n32983_o)
      n33021_q <= n33018_o;
    else
      n33021_q <= n33016_o;
endmodule

module delayi_2_8
  (input  clock_in,
   input  reset_in,
   input  [1:0] in_in,
   input  enable_in,
   output [1:0] out_out);
  wire [15:0] fifo_r;
  wire [1:0] n32937_o;
  wire n32940_o;
  wire [1:0] n32950_o;
  wire [1:0] n32951_o;
  wire [1:0] n32952_o;
  wire [1:0] n32953_o;
  wire [1:0] n32954_o;
  wire [1:0] n32955_o;
  wire [1:0] n32956_o;
  wire [1:0] n32957_o;
  wire [1:0] n32958_o;
  wire [1:0] n32959_o;
  wire [1:0] n32960_o;
  wire [1:0] n32961_o;
  wire [1:0] n32962_o;
  wire [1:0] n32963_o;
  wire [1:0] n32964_o;
  wire [1:0] n32965_o;
  wire [1:0] n32966_o;
  wire [1:0] n32967_o;
  wire [1:0] n32968_o;
  wire [1:0] n32969_o;
  wire [1:0] n32970_o;
  wire [1:0] n32971_o;
  wire [1:0] n32972_o;
  wire [15:0] n32973_o;
  wire [15:0] n32975_o;
  reg [15:0] n32978_q;
  assign out_out = n32937_o;
  /* ../../HW/src/util/delayi.vhd:46:8  */
  assign fifo_r = n32978_q; // (signal)
  /* ../../HW/src/util/delayi.vhd:48:18  */
  assign n32937_o = fifo_r[1:0];
  /* ../../HW/src/util/delayi.vhd:51:16  */
  assign n32940_o = ~reset_in;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32950_o = fifo_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32951_o = fifo_r[1:0];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32952_o = enable_in ? n32950_o : n32951_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32953_o = fifo_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32954_o = fifo_r[3:2];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32955_o = enable_in ? n32953_o : n32954_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32956_o = fifo_r[7:6];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32957_o = fifo_r[5:4];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32958_o = enable_in ? n32956_o : n32957_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32959_o = fifo_r[9:8];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32960_o = fifo_r[7:6];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32961_o = enable_in ? n32959_o : n32960_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32962_o = fifo_r[11:10];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32963_o = fifo_r[9:8];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32964_o = enable_in ? n32962_o : n32963_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32965_o = fifo_r[13:12];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32966_o = fifo_r[11:10];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32967_o = enable_in ? n32965_o : n32966_o;
  /* ../../HW/src/util/delayi.vhd:60:44  */
  assign n32968_o = fifo_r[15:14];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32969_o = fifo_r[13:12];
  /* ../../HW/src/util/delayi.vhd:59:21  */
  assign n32970_o = enable_in ? n32968_o : n32969_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32971_o = fifo_r[15:14];
  /* ../../HW/src/util/delayi.vhd:64:13  */
  assign n32972_o = enable_in ? in_in : n32971_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32973_o = {n32972_o, n32970_o, n32967_o, n32964_o, n32961_o, n32958_o, n32955_o, n32952_o};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32975_o = {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00};
  /* ../../HW/src/util/delayi.vhd:56:9  */
  always @(posedge clock_in or posedge n32940_o)
    if (n32940_o)
      n32978_q <= n32975_o;
    else
      n32978_q <= n32973_o;
endmodule

module delay_8
  (input  clock_in,
   input  reset_in,
   input  in_in,
   input  enable_in,
   output out_out);
  wire [7:0] fifo_r;
  wire n32894_o;
  wire n32897_o;
  wire n32907_o;
  wire n32908_o;
  wire n32909_o;
  wire n32910_o;
  wire n32911_o;
  wire n32912_o;
  wire n32913_o;
  wire n32914_o;
  wire n32915_o;
  wire n32916_o;
  wire n32917_o;
  wire n32918_o;
  wire n32919_o;
  wire n32920_o;
  wire n32921_o;
  wire n32922_o;
  wire n32923_o;
  wire n32924_o;
  wire n32925_o;
  wire n32926_o;
  wire n32927_o;
  wire n32928_o;
  wire n32929_o;
  wire [7:0] n32930_o;
  wire [7:0] n32932_o;
  reg [7:0] n32935_q;
  assign out_out = n32894_o;
  /* ../../HW/src/util/delay.vhd:46:8  */
  assign fifo_r = n32935_q; // (signal)
  /* ../../HW/src/util/delay.vhd:48:18  */
  assign n32894_o = fifo_r[0];
  /* ../../HW/src/util/delay.vhd:51:16  */
  assign n32897_o = ~reset_in;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32907_o = fifo_r[1];
  /* ../../HW/src/dp/dp_gen.vhd:776:5  */
  assign n32908_o = fifo_r[0];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32909_o = enable_in ? n32907_o : n32908_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32910_o = fifo_r[2];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32911_o = fifo_r[1];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32912_o = enable_in ? n32910_o : n32911_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32913_o = fifo_r[3];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32914_o = fifo_r[2];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32915_o = enable_in ? n32913_o : n32914_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32916_o = fifo_r[4];
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32917_o = fifo_r[3];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32918_o = enable_in ? n32916_o : n32917_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32919_o = fifo_r[5];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32920_o = fifo_r[4];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32921_o = enable_in ? n32919_o : n32920_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32922_o = fifo_r[6];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32923_o = fifo_r[5];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32924_o = enable_in ? n32922_o : n32923_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n32925_o = fifo_r[7];
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32926_o = fifo_r[6];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n32927_o = enable_in ? n32925_o : n32926_o;
  assign n32928_o = fifo_r[7];
  /* ../../HW/src/util/delay.vhd:64:13  */
  assign n32929_o = enable_in ? in_in : n32928_o;
  assign n32930_o = {n32929_o, n32927_o, n32924_o, n32921_o, n32918_o, n32915_o, n32912_o, n32909_o};
  assign n32932_o = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  /* ../../HW/src/util/delay.vhd:56:9  */
  always @(posedge clock_in or posedge n32897_o)
    if (n32897_o)
      n32935_q <= n32932_o;
    else
      n32935_q <= n32930_o;
endmodule

module dp_gen_3_1_5b55ec37559bb110228a6591713076b7fa2ce5e8
  (input  clock_in,
   input  reset_in,
   input  instruction_valid_in,
   input  instruction_latch_in,
   input  [23:0] instruction_source_in_stride0,
   input  [23:0] instruction_source_in_stride0_count,
   input  [24:0] instruction_source_in_stride0_max,
   input  [24:0] instruction_source_in_stride0_min,
   input  [23:0] instruction_source_in_stride1,
   input  [23:0] instruction_source_in_stride1_count,
   input  [24:0] instruction_source_in_stride1_max,
   input  [24:0] instruction_source_in_stride1_min,
   input  [23:0] instruction_source_in_stride2,
   input  [23:0] instruction_source_in_stride2_count,
   input  [24:0] instruction_source_in_stride2_max,
   input  [24:0] instruction_source_in_stride2_min,
   input  [23:0] instruction_source_in_stride3,
   input  [23:0] instruction_source_in_stride3_count,
   input  [24:0] instruction_source_in_stride3_max,
   input  [24:0] instruction_source_in_stride3_min,
   input  [23:0] instruction_source_in_stride4,
   input  [23:0] instruction_source_in_stride4_count,
   input  [24:0] instruction_source_in_stride4_max,
   input  [24:0] instruction_source_in_stride4_min,
   input  [24:0] instruction_source_in_burst_max,
   input  [24:0] instruction_source_in_burst_max2,
   input  [24:0] instruction_source_in_burst_max_init,
   input  [2:0] instruction_source_in_burst_max_index,
   input  [24:0] instruction_source_in_burst_min,
   input  [31:0] instruction_source_in_bar,
   input  [23:0] instruction_source_in_count,
   input  [23:0] instruction_source_in_burststride,
   input  instruction_source_in_double_precision,
   input  [1:0] instruction_source_in_data_model,
   input  instruction_source_in_scatter,
   input  [23:0] instruction_source_in_totalcount,
   input  [5:0] instruction_source_in_mcast,
   input  [15:0] instruction_source_in_data,
   input  instruction_source_in_repeat,
   input  [1:0] instruction_source_in_datatype,
   input  [1:0] instruction_source_in_bus_id,
   input  [23:0] instruction_source_in_bufsize,
   input  [23:0] instruction_source_in_burst_max_len,
   input  [23:0] instruction_dest_in_stride0,
   input  [23:0] instruction_dest_in_stride0_count,
   input  [24:0] instruction_dest_in_stride0_max,
   input  [24:0] instruction_dest_in_stride0_min,
   input  [23:0] instruction_dest_in_stride1,
   input  [23:0] instruction_dest_in_stride1_count,
   input  [24:0] instruction_dest_in_stride1_max,
   input  [24:0] instruction_dest_in_stride1_min,
   input  [23:0] instruction_dest_in_stride2,
   input  [23:0] instruction_dest_in_stride2_count,
   input  [24:0] instruction_dest_in_stride2_max,
   input  [24:0] instruction_dest_in_stride2_min,
   input  [23:0] instruction_dest_in_stride3,
   input  [23:0] instruction_dest_in_stride3_count,
   input  [24:0] instruction_dest_in_stride3_max,
   input  [24:0] instruction_dest_in_stride3_min,
   input  [23:0] instruction_dest_in_stride4,
   input  [23:0] instruction_dest_in_stride4_count,
   input  [24:0] instruction_dest_in_stride4_max,
   input  [24:0] instruction_dest_in_stride4_min,
   input  [24:0] instruction_dest_in_burst_max,
   input  [24:0] instruction_dest_in_burst_max2,
   input  [24:0] instruction_dest_in_burst_max_init,
   input  [2:0] instruction_dest_in_burst_max_index,
   input  [24:0] instruction_dest_in_burst_min,
   input  [31:0] instruction_dest_in_bar,
   input  [23:0] instruction_dest_in_count,
   input  [23:0] instruction_dest_in_burststride,
   input  instruction_dest_in_double_precision,
   input  [1:0] instruction_dest_in_data_model,
   input  instruction_dest_in_scatter,
   input  [23:0] instruction_dest_in_totalcount,
   input  [5:0] instruction_dest_in_mcast,
   input  [15:0] instruction_dest_in_data,
   input  instruction_dest_in_repeat,
   input  [1:0] instruction_dest_in_datatype,
   input  [1:0] instruction_dest_in_bus_id,
   input  [23:0] instruction_dest_in_bufsize,
   input  [23:0] instruction_dest_in_burst_max_len,
   input  instruction_stream_process_in,
   input  [1:0] instruction_stream_process_id_in,
   input  instruction_vm_in,
   input  [23:0] pre_instruction_source_in_stride0,
   input  [23:0] pre_instruction_source_in_stride0_count,
   input  [24:0] pre_instruction_source_in_stride0_max,
   input  [24:0] pre_instruction_source_in_stride0_min,
   input  [23:0] pre_instruction_source_in_stride1,
   input  [23:0] pre_instruction_source_in_stride1_count,
   input  [24:0] pre_instruction_source_in_stride1_max,
   input  [24:0] pre_instruction_source_in_stride1_min,
   input  [23:0] pre_instruction_source_in_stride2,
   input  [23:0] pre_instruction_source_in_stride2_count,
   input  [24:0] pre_instruction_source_in_stride2_max,
   input  [24:0] pre_instruction_source_in_stride2_min,
   input  [23:0] pre_instruction_source_in_stride3,
   input  [23:0] pre_instruction_source_in_stride3_count,
   input  [24:0] pre_instruction_source_in_stride3_max,
   input  [24:0] pre_instruction_source_in_stride3_min,
   input  [23:0] pre_instruction_source_in_stride4,
   input  [23:0] pre_instruction_source_in_stride4_count,
   input  [24:0] pre_instruction_source_in_stride4_max,
   input  [24:0] pre_instruction_source_in_stride4_min,
   input  [24:0] pre_instruction_source_in_burst_max,
   input  [24:0] pre_instruction_source_in_burst_max2,
   input  [24:0] pre_instruction_source_in_burst_max_init,
   input  [2:0] pre_instruction_source_in_burst_max_index,
   input  [24:0] pre_instruction_source_in_burst_min,
   input  [31:0] pre_instruction_source_in_bar,
   input  [23:0] pre_instruction_source_in_count,
   input  [23:0] pre_instruction_source_in_burststride,
   input  pre_instruction_source_in_double_precision,
   input  [1:0] pre_instruction_source_in_data_model,
   input  pre_instruction_source_in_scatter,
   input  [23:0] pre_instruction_source_in_totalcount,
   input  [5:0] pre_instruction_source_in_mcast,
   input  [15:0] pre_instruction_source_in_data,
   input  pre_instruction_source_in_repeat,
   input  [1:0] pre_instruction_source_in_datatype,
   input  [1:0] pre_instruction_source_in_bus_id,
   input  [23:0] pre_instruction_source_in_bufsize,
   input  [23:0] pre_instruction_source_in_burst_max_len,
   input  [23:0] pre_instruction_dest_in_stride0,
   input  [23:0] pre_instruction_dest_in_stride0_count,
   input  [24:0] pre_instruction_dest_in_stride0_max,
   input  [24:0] pre_instruction_dest_in_stride0_min,
   input  [23:0] pre_instruction_dest_in_stride1,
   input  [23:0] pre_instruction_dest_in_stride1_count,
   input  [24:0] pre_instruction_dest_in_stride1_max,
   input  [24:0] pre_instruction_dest_in_stride1_min,
   input  [23:0] pre_instruction_dest_in_stride2,
   input  [23:0] pre_instruction_dest_in_stride2_count,
   input  [24:0] pre_instruction_dest_in_stride2_max,
   input  [24:0] pre_instruction_dest_in_stride2_min,
   input  [23:0] pre_instruction_dest_in_stride3,
   input  [23:0] pre_instruction_dest_in_stride3_count,
   input  [24:0] pre_instruction_dest_in_stride3_max,
   input  [24:0] pre_instruction_dest_in_stride3_min,
   input  [23:0] pre_instruction_dest_in_stride4,
   input  [23:0] pre_instruction_dest_in_stride4_count,
   input  [24:0] pre_instruction_dest_in_stride4_max,
   input  [24:0] pre_instruction_dest_in_stride4_min,
   input  [24:0] pre_instruction_dest_in_burst_max,
   input  [24:0] pre_instruction_dest_in_burst_max2,
   input  [24:0] pre_instruction_dest_in_burst_max_init,
   input  [2:0] pre_instruction_dest_in_burst_max_index,
   input  [24:0] pre_instruction_dest_in_burst_min,
   input  [31:0] pre_instruction_dest_in_bar,
   input  [23:0] pre_instruction_dest_in_count,
   input  [23:0] pre_instruction_dest_in_burststride,
   input  pre_instruction_dest_in_double_precision,
   input  [1:0] pre_instruction_dest_in_data_model,
   input  pre_instruction_dest_in_scatter,
   input  [23:0] pre_instruction_dest_in_totalcount,
   input  [5:0] pre_instruction_dest_in_mcast,
   input  [15:0] pre_instruction_dest_in_data,
   input  pre_instruction_dest_in_repeat,
   input  [1:0] pre_instruction_dest_in_datatype,
   input  [1:0] pre_instruction_dest_in_bus_id,
   input  [23:0] pre_instruction_dest_in_bufsize,
   input  [23:0] pre_instruction_dest_in_burst_max_len,
   input  [1:0] pre_instruction_bus_id_source_in,
   input  [1:0] pre_instruction_bus_id_dest_in,
   input  instruction_source_addr_mode_in,
   input  instruction_dest_addr_mode_in,
   input  [1:0] instruction_bus_id_source_in,
   input  [1:0] instruction_data_type_source_in,
   input  [1:0] instruction_data_model_source_in,
   input  [1:0] instruction_bus_id_dest_in,
   input  [1:0] instruction_data_type_dest_in,
   input  [1:0] instruction_data_model_dest_in,
   input  [23:0] instruction_gen_len_in,
   input  [5:0] instruction_mcast_in,
   input  instruction_thread_in,
   input  [15:0] instruction_data_in,
   input  instruction_repeat_in,
   input  [14:0] wr_maxburstlen_in,
   input  [2:0] wr_full_in,
   input  [2:0] waitreq_in,
   input  [71:0] gen_bar_in,
   output ready_out,
   output [2:0] gen_valid_out,
   output gen_vm_out,
   output gen_fork_out,
   output [1:0] gen_data_flow_out,
   output gen_src_stream_out,
   output gen_dest_stream_out,
   output [1:0] gen_stream_id_out,
   output [2:0] gen_src_vector_out,
   output [2:0] gen_dst_vector_out,
   output [1:0] gen_src_scatter_out,
   output [1:0] gen_dst_scatter_out,
   output [3:0] gen_src_start_out,
   output [3:0] gen_src_end_out,
   output [3:0] gen_dst_end_out,
   output [31:0] gen_addr_source_out,
   output gen_addr_source_mode_out,
   output [31:0] gen_addr_dest_out,
   output gen_addr_dest_mode_out,
   output gen_eof_out,
   output [1:0] gen_bus_id_source_out,
   output [1:0] gen_data_type_source_out,
   output [1:0] gen_data_model_source_out,
   output [1:0] gen_bus_id_dest_out,
   output gen_busy_dest_out,
   output [1:0] gen_data_type_dest_out,
   output [1:0] gen_data_model_dest_out,
   output [4:0] gen_burstlen_source_out,
   output [4:0] gen_burstlen_dest_out,
   output gen_thread_out,
   output [5:0] gen_mcast_out,
   output [63:0] gen_data_out,
   output [31:0] log_out,
   output log_valid_out);
  wire [775:0] n29602_o;
  wire [775:0] n29603_o;
  wire [775:0] n29604_o;
  wire [775:0] n29605_o;
  wire [775:0] s_template_r;
  wire [23:0] s_i0_r;
  wire [23:0] s_i1_r;
  wire [23:0] s_i2_r;
  wire [23:0] s_i3_r;
  wire [23:0] s_i4_r;
  wire [23:0] s_i0_count_r;
  wire [23:0] s_i1_count_r;
  wire [23:0] s_i2_count_r;
  wire [23:0] s_i3_count_r;
  wire [23:0] s_i4_count_r;
  wire [23:0] s_burstlen_r;
  wire [23:0] s_burstpos_r;
  reg [23:0] s_burstremain_r;
  reg s_valid_r;
  wire [24:0] s_i0_start_r;
  wire [24:0] s_i1_start_r;
  wire [24:0] s_i2_start_r;
  wire [24:0] s_i3_start_r;
  wire [24:0] s_i4_start_r;
  wire [23:0] s_burstpos_stride_r;
  wire [24:0] s_burstpos_start_r;
  wire [3:0] s_burstpos_start_rr;
  wire [3:0] s_burstpos_start_rrr;
  wire [3:0] s_burstpos_start_rrrr;
  wire [26:0] s_burstpos_end_r;
  wire [3:0] s_burstpos_end_rr;
  wire [3:0] s_burstpos_end_rrr;
  wire [26:0] d_burstpos_end_r;
  wire [3:0] d_burstpos_end_rr;
  wire [3:0] d_burstpos_end_rrr;
  wire [775:0] d_template_r;
  wire [23:0] d_i0_r;
  wire [23:0] d_i1_r;
  wire [23:0] d_i2_r;
  wire [23:0] d_i3_r;
  wire [23:0] d_i4_r;
  wire [23:0] d_i0_count_r;
  wire [23:0] d_i1_count_r;
  wire [23:0] d_i2_count_r;
  wire [23:0] d_i3_count_r;
  wire [23:0] d_i4_count_r;
  wire [24:0] d_burst_max_r;
  wire [23:0] d_burstlen_r;
  wire [23:0] d_burstpos_r;
  reg [23:0] d_burstremain_r;
  reg d_valid_r;
  wire [23:0] currlen_r;
  wire [23:0] currlen_new;
  wire reload;
  wire s_burstlen_wrap;
  wire s_i0_wrap;
  wire s_i1_wrap;
  wire s_i2_wrap;
  wire s_i3_wrap;
  wire s_i4_wrap;
  wire [23:0] s_burstlen_new;
  wire [23:0] s_burstpos_new;
  wire [23:0] s_i0_new;
  wire [23:0] s_i1_new;
  wire [23:0] s_i2_new;
  wire [23:0] s_i3_new;
  wire [23:0] s_i4_new;
  wire [23:0] s_i0_count_new;
  wire [23:0] s_i1_count_new;
  wire [23:0] s_i2_count_new;
  wire [23:0] s_i3_count_new;
  wire [23:0] s_i4_count_new;
  wire [24:0] s_burstpos_start_new;
  wire [24:0] s_i0_start_new;
  wire [24:0] s_i1_start_new;
  wire [24:0] s_i2_start_new;
  wire [24:0] s_i3_start_new;
  wire [24:0] s_i4_start_new;
  wire d_burstlen_wrap;
  wire d_i0_wrap;
  wire d_i1_wrap;
  wire d_i2_wrap;
  wire d_i3_wrap;
  wire d_i4_wrap;
  wire [23:0] d_burstlen_new;
  wire [23:0] d_burstpos_new;
  wire [23:0] d_i0_new;
  wire [23:0] d_i1_new;
  wire [23:0] d_i2_new;
  wire [23:0] d_i3_new;
  wire [23:0] d_i4_new;
  wire [23:0] d_i0_new2;
  wire [23:0] d_i1_new2;
  wire [23:0] d_i2_new2;
  wire [23:0] d_i3_new2;
  wire [23:0] d_i4_new2;
  wire [23:0] d_i0_count_new;
  wire [23:0] d_i1_count_new;
  wire [23:0] d_i2_count_new;
  wire [23:0] d_i3_count_new;
  wire [23:0] d_i4_count_new;
  wire running_r;
  wire running_rr;
  wire running_rrr;
  wire running_rrrr;
  wire [2:0] gen_valid_r;
  wire [1:0] dp_dst_bus_id_r;
  wire [1:0] dp_dst_bus_id_rr;
  wire [1:0] dp_dst_bus_id_rrr;
  wire [1:0] dp_dst_bus_id_rrrr;
  wire [1:0] dp_src_bus_id_r;
  wire [1:0] dp_src_bus_id_rr;
  wire [1:0] dp_src_bus_id_rrr;
  wire [1:0] dp_src_bus_id_rrrr;
  wire [1:0] dp_dst_data_type_r;
  wire [1:0] dp_dst_data_type_rr;
  wire [1:0] dp_dst_data_type_rrr;
  wire [1:0] dp_dst_data_type_rrrr;
  wire [1:0] dp_src_data_type_r;
  wire [1:0] dp_src_data_type_rr;
  wire [1:0] dp_src_data_type_rrr;
  wire [1:0] dp_src_data_type_rrrr;
  wire [1:0] dp_src_data_model_r;
  wire [1:0] dp_src_data_model_rr;
  wire [1:0] dp_src_data_model_rrr;
  wire [1:0] dp_src_data_model_rrrr;
  wire [1:0] dp_dst_data_model_r;
  wire [1:0] dp_dst_data_model_rr;
  wire [1:0] dp_dst_data_model_rrr;
  wire [1:0] dp_dst_data_model_rrrr;
  wire dp_thread_r;
  wire dp_thread_rr;
  wire dp_thread_rrr;
  wire dp_thread_rrrr;
  reg [5:0] dp_mcast_r;
  reg [5:0] dp_mcast_rr;
  reg [5:0] dp_mcast_rrr;
  reg [5:0] dp_mcast_rrrr;
  wire [63:0] data_r;
  wire [63:0] data_rr;
  wire [63:0] data_rrr;
  wire [63:0] data_rrrr;
  wire [23:0] s_bufsize_r;
  wire [23:0] s_bufsize_rr;
  wire [23:0] s_temp1_r;
  wire [31:0] s_temp2_r;
  wire [23:0] s_temp3_r;
  wire [23:0] s_temp4_r;
  wire [23:0] s_temp5_r;
  wire [31:0] s_temp4_rr;
  wire [31:0] s_gen_addr_r;
  wire [4:0] s_gen_burstlen_r;
  wire [4:0] s_gen_burstlen_rr;
  wire s_gen_burstlen_progress_r;
  wire s_i0_valid;
  wire s_i1_valid;
  wire s_i2_valid;
  wire s_i3_valid;
  wire s_i4_valid;
  wire s_burst_valid;
  wire s_i0_start_valid;
  wire s_i1_start_valid;
  wire s_i2_start_valid;
  wire s_i3_start_valid;
  wire s_i4_start_valid;
  wire s_burst_start_valid;
  wire [23:0] d_bufsize_r;
  wire [23:0] d_bufsize_rr;
  wire [23:0] d_temp1_r;
  wire [31:0] d_temp2_r;
  wire [23:0] d_temp3_r;
  wire [23:0] d_temp4_r;
  wire [23:0] d_temp5_r;
  wire [31:0] d_temp4_rr;
  wire [31:0] d_gen_addr_r;
  wire [4:0] d_gen_burstlen_r;
  wire [4:0] d_gen_burstlen_rr;
  wire d_i0_valid;
  wire d_i1_valid;
  wire d_i2_valid;
  wire d_i3_valid;
  wire d_i4_valid;
  wire d_burst_valid;
  wire eof_r;
  wire eof_rr;
  wire eof_rrr;
  wire eof_rrrr;
  reg done_r;
  wire repeat_r;
  wire [1:0] data_flow_r;
  wire [1:0] data_flow_rr;
  wire [1:0] data_flow_rrr;
  wire [1:0] data_flow_rrrr;
  wire stream_src_r;
  wire stream_src_rr;
  wire stream_src_rrr;
  wire stream_src_rrrr;
  wire stream_dest_r;
  wire stream_dest_rr;
  wire stream_dest_rrr;
  wire stream_dest_rrrr;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire [1:0] stream_id_r;
  wire [1:0] stream_id_rr;
  wire [1:0] stream_id_rrr;
  wire [1:0] stream_id_rrrr;
  wire src_double_r;
  wire src_double_rr;
  wire src_double_rrr;
  wire dst_double_r;
  wire dst_double_rr;
  wire dst_double_rrr;
  wire [2:0] src_vector_r;
  wire [2:0] src_vector_rr;
  wire [2:0] src_vector_rrr;
  wire [2:0] src_vector_rrrr;
  wire [2:0] dst_vector_r;
  wire [2:0] dst_vector_rr;
  wire [2:0] dst_vector_rrr;
  wire [2:0] dst_vector_rrrr;
  wire src_addr_mode_r;
  wire src_addr_mode_rr;
  wire src_addr_mode_rrr;
  wire src_addr_mode_rrrr;
  wire dst_addr_mode_r;
  wire dst_addr_mode_rr;
  wire dst_addr_mode_rrr;
  wire dst_addr_mode_rrrr;
  wire [1:0] src_scatter_r;
  wire [1:0] src_scatter_rr;
  wire [1:0] src_scatter_rrr;
  wire [1:0] src_scatter_rrrr;
  wire [1:0] dst_scatter_r;
  wire [1:0] dst_scatter_rr;
  wire [1:0] dst_scatter_rrr;
  wire [1:0] dst_scatter_rrrr;
  wire [2:0] src_vector;
  wire [2:0] dst_vector;
  wire [1:0] src_scatter;
  wire [1:0] dst_scatter;
  wire src_is_burst_r;
  wire src_is_burst_rr;
  wire dst_is_burst_r;
  wire dst_is_burst_rr;
  wire [2:0] src_is_vector_r;
  wire [2:0] dst_is_vector_r;
  wire [5:0] src_is_scatter_r;
  wire [5:0] dst_is_scatter_r;
  wire [24:0] s_burst_actual_max_r;
  wire [31:0] log;
  wire [31:0] log_r;
  wire log_valid_r;
  wire source_double_precision;
  wire dest_double_precision;
  wire waitreq;
  wire ready;
  wire gen_busy_dest_r;
  wire n29648_o;
  wire n29650_o;
  wire n29651_o;
  wire n29653_o;
  wire n29655_o;
  wire n29656_o;
  wire n29659_o;
  wire n29660_o;
  wire n29661_o;
  wire n29662_o;
  wire n29663_o;
  wire n29664_o;
  wire n29665_o;
  wire n29666_o;
  wire n29667_o;
  wire n29670_o;
  wire n29671_o;
  wire n29672_o;
  wire [23:0] n29675_o;
  wire n29686_o;
  wire [2:0] n29688_o;
  wire n29690_o;
  wire n29692_o;
  wire n29693_o;
  wire n29694_o;
  wire n29695_o;
  wire [23:0] n29696_o;
  wire n29698_o;
  wire [23:0] n29700_o;
  wire n29702_o;
  wire [1:0] n29705_o;
  wire [1:0] n29706_o;
  wire [1:0] n29707_o;
  wire [2:0] n29708_o;
  wire n29710_o;
  wire n29712_o;
  wire n29713_o;
  wire n29714_o;
  wire n29715_o;
  wire [23:0] n29716_o;
  wire n29718_o;
  wire [23:0] n29719_o;
  wire n29721_o;
  wire [1:0] n29722_o;
  wire [1:0] n29723_o;
  wire [1:0] n29724_o;
  wire n29726_o;
  wire [23:0] n29727_o;
  wire n29729_o;
  wire [23:0] n29730_o;
  wire n29732_o;
  wire [2:0] n29733_o;
  wire n29735_o;
  wire n29736_o;
  wire n29737_o;
  wire n29740_o;
  wire [23:0] n29741_o;
  wire n29743_o;
  wire [2:0] n29744_o;
  wire n29746_o;
  wire [2:0] n29747_o;
  wire n29749_o;
  wire n29750_o;
  wire [2:0] n29751_o;
  wire n29753_o;
  wire n29754_o;
  wire [2:0] n29755_o;
  wire n29757_o;
  wire n29758_o;
  wire [2:0] n29759_o;
  wire n29761_o;
  wire n29762_o;
  wire [23:0] n29763_o;
  wire n29765_o;
  wire n29766_o;
  wire [2:0] n29767_o;
  wire n29769_o;
  wire n29770_o;
  wire [2:0] n29771_o;
  wire n29773_o;
  wire n29774_o;
  wire [2:0] n29775_o;
  wire n29777_o;
  wire n29778_o;
  wire n29779_o;
  wire n29782_o;
  wire n29783_o;
  wire n29785_o;
  wire [23:0] n29786_o;
  wire n29788_o;
  wire [23:0] n29789_o;
  wire n29791_o;
  wire [2:0] n29792_o;
  wire n29794_o;
  wire n29795_o;
  wire n29796_o;
  wire n29799_o;
  wire [23:0] n29800_o;
  wire n29802_o;
  wire [2:0] n29803_o;
  wire n29805_o;
  wire [2:0] n29806_o;
  wire n29808_o;
  wire n29809_o;
  wire [2:0] n29810_o;
  wire n29812_o;
  wire n29813_o;
  wire [2:0] n29814_o;
  wire n29816_o;
  wire n29817_o;
  wire [2:0] n29818_o;
  wire n29820_o;
  wire n29821_o;
  wire [23:0] n29822_o;
  wire n29824_o;
  wire n29825_o;
  wire [2:0] n29826_o;
  wire n29828_o;
  wire n29829_o;
  wire [2:0] n29830_o;
  wire n29832_o;
  wire n29833_o;
  wire [2:0] n29834_o;
  wire n29836_o;
  wire n29837_o;
  wire n29838_o;
  wire n29841_o;
  wire n29842_o;
  wire [1:0] n29843_o;
  wire n29845_o;
  wire n29847_o;
  wire n29848_o;
  wire n29849_o;
  wire n29850_o;
  wire [23:0] n29851_o;
  wire n29853_o;
  wire [23:0] n29854_o;
  wire n29856_o;
  wire [1:0] n29857_o;
  wire [1:0] n29858_o;
  wire [1:0] n29859_o;
  wire [1:0] n29860_o;
  wire n29862_o;
  wire n29864_o;
  wire n29865_o;
  wire n29866_o;
  wire n29867_o;
  wire [23:0] n29868_o;
  wire n29870_o;
  wire [23:0] n29871_o;
  wire n29873_o;
  wire [1:0] n29874_o;
  wire [1:0] n29875_o;
  wire [1:0] n29876_o;
  wire n29878_o;
  wire [23:0] n29879_o;
  wire n29881_o;
  wire [23:0] n29882_o;
  wire n29884_o;
  wire [1:0] n29885_o;
  wire n29887_o;
  wire n29888_o;
  wire n29889_o;
  wire n29892_o;
  wire [23:0] n29893_o;
  wire n29895_o;
  wire [1:0] n29896_o;
  wire n29898_o;
  wire [1:0] n29899_o;
  wire n29901_o;
  wire n29902_o;
  wire [1:0] n29903_o;
  wire n29905_o;
  wire n29906_o;
  wire [1:0] n29907_o;
  wire n29909_o;
  wire n29910_o;
  wire [1:0] n29911_o;
  wire n29913_o;
  wire n29914_o;
  wire [23:0] n29915_o;
  wire n29917_o;
  wire n29918_o;
  wire [1:0] n29919_o;
  wire n29921_o;
  wire n29922_o;
  wire [1:0] n29923_o;
  wire n29925_o;
  wire n29926_o;
  wire [1:0] n29927_o;
  wire n29929_o;
  wire n29930_o;
  wire n29931_o;
  wire n29934_o;
  wire n29935_o;
  wire n29937_o;
  wire [23:0] n29938_o;
  wire n29940_o;
  wire [23:0] n29941_o;
  wire n29943_o;
  wire [1:0] n29944_o;
  wire n29946_o;
  wire n29947_o;
  wire n29948_o;
  wire n29951_o;
  wire [23:0] n29952_o;
  wire n29954_o;
  wire [1:0] n29955_o;
  wire n29957_o;
  wire [1:0] n29958_o;
  wire n29960_o;
  wire n29961_o;
  wire [1:0] n29962_o;
  wire n29964_o;
  wire n29965_o;
  wire [1:0] n29966_o;
  wire n29968_o;
  wire n29969_o;
  wire [1:0] n29970_o;
  wire n29972_o;
  wire n29973_o;
  wire [23:0] n29974_o;
  wire n29976_o;
  wire n29977_o;
  wire [1:0] n29978_o;
  wire n29980_o;
  wire n29981_o;
  wire [1:0] n29982_o;
  wire n29984_o;
  wire n29985_o;
  wire [1:0] n29986_o;
  wire n29988_o;
  wire n29989_o;
  wire n29990_o;
  wire n29993_o;
  wire n29994_o;
  wire n29995_o;
  wire n29997_o;
  wire n29999_o;
  wire n30000_o;
  wire n30001_o;
  wire n30002_o;
  wire [23:0] n30003_o;
  wire n30005_o;
  wire [23:0] n30006_o;
  wire n30008_o;
  wire [1:0] n30009_o;
  wire [1:0] n30010_o;
  wire [1:0] n30011_o;
  wire n30012_o;
  wire n30014_o;
  wire n30016_o;
  wire n30017_o;
  wire n30018_o;
  wire n30019_o;
  wire [23:0] n30020_o;
  wire n30022_o;
  wire [23:0] n30023_o;
  wire n30025_o;
  wire [1:0] n30026_o;
  wire [1:0] n30027_o;
  wire [1:0] n30028_o;
  wire n30030_o;
  wire [23:0] n30031_o;
  wire n30033_o;
  wire [23:0] n30034_o;
  wire n30036_o;
  wire n30037_o;
  wire n30039_o;
  wire n30040_o;
  wire n30041_o;
  wire n30044_o;
  wire [23:0] n30045_o;
  wire n30047_o;
  wire n30048_o;
  wire n30050_o;
  wire n30051_o;
  wire n30053_o;
  wire n30054_o;
  wire n30055_o;
  wire n30057_o;
  wire n30058_o;
  wire n30059_o;
  wire n30061_o;
  wire n30062_o;
  wire n30063_o;
  wire n30065_o;
  wire n30066_o;
  wire [23:0] n30067_o;
  wire n30069_o;
  wire n30070_o;
  wire n30071_o;
  wire n30073_o;
  wire n30074_o;
  wire n30075_o;
  wire n30077_o;
  wire n30078_o;
  wire n30079_o;
  wire n30081_o;
  wire n30082_o;
  wire n30083_o;
  wire n30086_o;
  wire n30087_o;
  wire n30089_o;
  wire [23:0] n30090_o;
  wire n30092_o;
  wire [23:0] n30093_o;
  wire n30095_o;
  wire n30096_o;
  wire n30098_o;
  wire n30099_o;
  wire n30100_o;
  wire n30103_o;
  wire [23:0] n30104_o;
  wire n30106_o;
  wire n30107_o;
  wire n30109_o;
  wire n30110_o;
  wire n30112_o;
  wire n30113_o;
  wire n30114_o;
  wire n30116_o;
  wire n30117_o;
  wire n30118_o;
  wire n30120_o;
  wire n30121_o;
  wire n30122_o;
  wire n30124_o;
  wire n30125_o;
  wire [23:0] n30126_o;
  wire n30128_o;
  wire n30129_o;
  wire n30130_o;
  wire n30132_o;
  wire n30133_o;
  wire n30134_o;
  wire n30136_o;
  wire n30137_o;
  wire n30138_o;
  wire n30140_o;
  wire n30141_o;
  wire n30142_o;
  wire n30145_o;
  wire n30146_o;
  wire [2:0] n30147_o;
  wire [2:0] n30149_o;
  wire [5:0] n30151_o;
  wire [5:0] n30153_o;
  wire n30172_o;
  wire [1:0] n30173_o;
  wire n30175_o;
  wire n30176_o;
  wire n30177_o;
  wire n30178_o;
  wire n30179_o;
  wire n30180_o;
  wire [1:0] n30181_o;
  wire n30183_o;
  wire n30184_o;
  wire n30185_o;
  wire n30186_o;
  wire n30187_o;
  wire n30188_o;
  wire [1:0] n30189_o;
  wire [1:0] n30190_o;
  wire n30191_o;
  wire [1:0] n30192_o;
  wire n30194_o;
  wire n30195_o;
  wire n30196_o;
  wire [1:0] n30197_o;
  wire n30199_o;
  wire n30200_o;
  wire n30201_o;
  wire [1:0] n30202_o;
  wire [1:0] n30203_o;
  wire n30204_o;
  wire [1:0] n30205_o;
  wire n30207_o;
  wire n30208_o;
  wire n30209_o;
  wire [1:0] n30210_o;
  wire n30212_o;
  wire n30213_o;
  wire n30214_o;
  wire [1:0] n30215_o;
  wire [1:0] n30216_o;
  wire [2:0] n30219_o;
  wire [2:0] n30222_o;
  wire [1:0] n30224_o;
  wire [1:0] n30226_o;
  wire [2:0] n30228_o;
  wire [2:0] n30230_o;
  wire [1:0] n30231_o;
  wire [1:0] n30232_o;
  wire [2:0] n30234_o;
  wire [2:0] n30236_o;
  wire [1:0] n30237_o;
  wire [1:0] n30238_o;
  wire [23:0] n30241_o;
  wire [23:0] n30242_o;
  wire [23:0] n30243_o;
  wire [23:0] n30244_o;
  wire [23:0] n30245_o;
  wire [23:0] n30246_o;
  wire [23:0] n30247_o;
  wire [23:0] n30248_o;
  wire [23:0] n30249_o;
  wire [23:0] n30250_o;
  wire [23:0] n30251_o;
  wire [23:0] n30252_o;
  wire [23:0] n30253_o;
  wire [24:0] n30255_o;
  wire [24:0] n30256_o;
  wire [23:0] n30257_o;
  wire [24:0] n30259_o;
  wire [24:0] n30260_o;
  wire [23:0] n30261_o;
  wire [24:0] n30263_o;
  wire [24:0] n30264_o;
  wire [23:0] n30265_o;
  wire [24:0] n30267_o;
  wire [24:0] n30268_o;
  wire [23:0] n30269_o;
  wire [24:0] n30271_o;
  wire [24:0] n30272_o;
  wire [23:0] n30273_o;
  wire [24:0] n30275_o;
  wire [24:0] n30276_o;
  wire [23:0] n30278_o;
  wire [23:0] n30280_o;
  wire [23:0] n30282_o;
  wire [23:0] n30284_o;
  wire [23:0] n30286_o;
  wire [23:0] n30288_o;
  wire [23:0] n30289_o;
  wire [23:0] n30290_o;
  wire [23:0] n30291_o;
  wire [23:0] n30292_o;
  wire [23:0] n30293_o;
  wire [23:0] n30294_o;
  wire [23:0] n30295_o;
  wire [23:0] n30296_o;
  wire [23:0] n30297_o;
  wire [23:0] n30298_o;
  wire [23:0] n30299_o;
  wire [23:0] n30300_o;
  wire [22:0] n30301_o;
  wire [23:0] n30303_o;
  wire [23:0] n30304_o;
  wire [22:0] n30305_o;
  wire [23:0] n30307_o;
  wire [23:0] n30308_o;
  wire [22:0] n30309_o;
  wire [23:0] n30311_o;
  wire [23:0] n30312_o;
  wire [22:0] n30313_o;
  wire [23:0] n30315_o;
  wire [23:0] n30316_o;
  wire [22:0] n30317_o;
  wire [23:0] n30319_o;
  wire [23:0] n30320_o;
  wire [23:0] n30322_o;
  wire [23:0] n30324_o;
  wire [23:0] n30326_o;
  wire [23:0] n30328_o;
  wire [23:0] n30330_o;
  localparam n30331_o = 1'b0;
  wire n30333_o;
  wire n30334_o;
  wire n30335_o;
  wire [2:0] n30338_o;
  wire n30340_o;
  wire n30341_o;
  wire [23:0] n30344_o;
  wire n30345_o;
  wire n30346_o;
  wire [23:0] n30349_o;
  wire n30350_o;
  wire n30351_o;
  wire [23:0] n30354_o;
  wire n30355_o;
  wire n30356_o;
  wire [23:0] n30359_o;
  wire n30360_o;
  wire n30361_o;
  wire [23:0] n30364_o;
  wire n30365_o;
  wire n30366_o;
  wire [23:0] n30369_o;
  wire n30370_o;
  wire n30371_o;
  wire [23:0] n30374_o;
  wire n30375_o;
  wire n30376_o;
  wire n30377_o;
  wire n30378_o;
  wire n30379_o;
  wire [23:0] n30382_o;
  wire n30383_o;
  wire n30384_o;
  wire n30385_o;
  wire n30386_o;
  wire n30387_o;
  wire [23:0] n30390_o;
  wire n30391_o;
  wire n30392_o;
  wire n30393_o;
  wire n30394_o;
  wire n30395_o;
  wire [23:0] n30398_o;
  wire n30399_o;
  wire n30400_o;
  wire n30401_o;
  wire n30402_o;
  wire n30403_o;
  wire [23:0] n30406_o;
  wire n30407_o;
  wire n30408_o;
  wire n30409_o;
  wire n30410_o;
  wire n30411_o;
  wire [23:0] n30414_o;
  wire n30415_o;
  wire n30416_o;
  wire n30417_o;
  wire n30418_o;
  wire n30419_o;
  wire n30421_o;
  wire n30422_o;
  wire n30423_o;
  wire n30424_o;
  wire n30425_o;
  wire n30426_o;
  wire n30427_o;
  wire n30428_o;
  wire n30429_o;
  wire n30430_o;
  wire [24:0] n30432_o;
  wire [24:0] n30433_o;
  wire n30435_o;
  wire n30436_o;
  wire [23:0] n30439_o;
  wire n30440_o;
  wire n30441_o;
  wire [23:0] n30444_o;
  wire n30445_o;
  wire n30446_o;
  wire [23:0] n30449_o;
  wire n30450_o;
  wire n30451_o;
  wire [23:0] n30454_o;
  wire n30455_o;
  wire n30456_o;
  wire [23:0] n30459_o;
  wire n30460_o;
  wire n30461_o;
  wire [23:0] n30464_o;
  wire n30465_o;
  wire n30466_o;
  wire [23:0] n30469_o;
  wire n30470_o;
  wire n30471_o;
  wire n30472_o;
  wire n30473_o;
  wire n30474_o;
  wire [23:0] n30477_o;
  wire n30478_o;
  wire n30479_o;
  wire n30480_o;
  wire n30481_o;
  wire n30482_o;
  wire [23:0] n30485_o;
  wire n30486_o;
  wire n30487_o;
  wire n30488_o;
  wire n30489_o;
  wire n30490_o;
  wire [23:0] n30493_o;
  wire n30494_o;
  wire n30495_o;
  wire n30496_o;
  wire n30497_o;
  wire n30498_o;
  wire [23:0] n30501_o;
  wire n30502_o;
  wire n30503_o;
  wire n30504_o;
  wire n30505_o;
  wire n30506_o;
  wire [23:0] n30509_o;
  wire n30510_o;
  wire n30511_o;
  wire n30512_o;
  wire n30513_o;
  wire n30514_o;
  wire n30526_o;
  wire n30528_o;
  wire n30530_o;
  wire n30532_o;
  wire n30534_o;
  wire n30536_o;
  wire n30538_o;
  wire n30540_o;
  wire [23:0] n30544_o;
  wire [23:0] n30545_o;
  wire [23:0] n30546_o;
  wire [31:0] n30547_o;
  wire [23:0] n30548_o;
  wire [23:0] n30549_o;
  wire [23:0] n30550_o;
  wire [23:0] n30551_o;
  wire [23:0] n30552_o;
  wire [31:0] n30553_o;
  wire [31:0] n30554_o;
  wire [31:0] n30556_o;
  wire [31:0] n30557_o;
  wire n30561_o;
  wire [4:0] n30565_o;
  wire n30567_o;
  wire n30570_o;
  wire [26:0] n30571_o;
  wire [23:0] n30572_o;
  wire [26:0] n30573_o;
  wire [26:0] n30574_o;
  wire [26:0] n30576_o;
  wire [26:0] n30578_o;
  wire [26:0] n30579_o;
  wire n30580_o;
  wire [22:0] n30581_o;
  wire n30583_o;
  wire [3:0] n30584_o;
  wire [3:0] n30586_o;
  wire [3:0] n30588_o;
  wire [22:0] n30589_o;
  wire [24:0] n30590_o;
  wire [24:0] n30591_o;
  wire [24:0] n30592_o;
  wire [24:0] n30594_o;
  wire [24:0] n30595_o;
  wire n30597_o;
  wire [24:0] n30598_o;
  wire n30599_o;
  wire [3:0] n30600_o;
  wire [3:0] n30601_o;
  wire [3:0] n30603_o;
  wire [22:0] n30605_o;
  wire [23:0] n30607_o;
  wire [23:0] n30608_o;
  wire n30610_o;
  wire [22:0] n30611_o;
  wire n30614_o;
  wire [21:0] n30615_o;
  wire n30618_o;
  wire [20:0] n30619_o;
  wire [23:0] n30621_o;
  wire [23:0] n30622_o;
  wire [23:0] n30623_o;
  wire [23:0] n30624_o;
  wire [23:0] n30625_o;
  wire [23:0] n30626_o;
  wire n30627_o;
  wire n30628_o;
  wire n30629_o;
  wire n30630_o;
  wire n30631_o;
  wire n30632_o;
  wire n30633_o;
  wire n30634_o;
  wire n30635_o;
  wire n30636_o;
  wire n30637_o;
  wire n30638_o;
  wire n30640_o;
  wire [18:0] n30641_o;
  wire n30643_o;
  wire [4:0] n30644_o;
  wire n30646_o;
  wire n30647_o;
  wire [4:0] n30648_o;
  wire [4:0] n30650_o;
  wire n30651_o;
  wire [18:0] n30652_o;
  wire n30654_o;
  wire [4:0] n30655_o;
  wire n30656_o;
  wire n30657_o;
  wire [4:0] n30658_o;
  wire [4:0] n30660_o;
  wire [4:0] n30662_o;
  wire [4:0] n30663_o;
  wire [4:0] n30665_o;
  wire n30666_o;
  wire [4:0] n30669_o;
  wire [4:0] n30670_o;
  wire [4:0] n30673_o;
  wire [1:0] n30675_o;
  wire [2:0] n30677_o;
  wire [2:0] n30678_o;
  wire n30679_o;
  wire n30680_o;
  wire [21:0] n30681_o;
  wire n30683_o;
  wire [3:0] n30684_o;
  wire [3:0] n30687_o;
  wire [3:0] n30688_o;
  wire [3:0] n30690_o;
  wire [1:0] n30691_o;
  wire [2:0] n30693_o;
  wire [2:0] n30694_o;
  wire [23:0] n30695_o;
  wire [23:0] n30696_o;
  wire [23:0] n30697_o;
  wire [31:0] n30698_o;
  wire [23:0] n30699_o;
  wire [23:0] n30700_o;
  wire [23:0] n30701_o;
  wire [23:0] n30702_o;
  wire [23:0] n30703_o;
  wire [31:0] n30704_o;
  wire [31:0] n30705_o;
  wire [31:0] n30707_o;
  wire [31:0] n30708_o;
  wire [26:0] n30709_o;
  wire [23:0] n30710_o;
  wire [26:0] n30711_o;
  wire [26:0] n30712_o;
  wire [26:0] n30714_o;
  wire [26:0] n30716_o;
  wire [26:0] n30717_o;
  wire n30718_o;
  wire [22:0] n30719_o;
  wire n30721_o;
  wire [3:0] n30722_o;
  wire [3:0] n30724_o;
  wire [3:0] n30726_o;
  wire [22:0] n30727_o;
  wire [24:0] n30728_o;
  wire [24:0] n30729_o;
  wire [24:0] n30730_o;
  wire [24:0] n30732_o;
  wire [24:0] n30733_o;
  wire n30735_o;
  wire [24:0] n30736_o;
  wire n30737_o;
  wire [3:0] n30738_o;
  wire [3:0] n30739_o;
  wire [3:0] n30741_o;
  wire [22:0] n30743_o;
  wire [23:0] n30745_o;
  wire [23:0] n30746_o;
  wire n30748_o;
  wire [22:0] n30749_o;
  wire n30752_o;
  wire [21:0] n30753_o;
  wire n30756_o;
  wire [20:0] n30757_o;
  wire [23:0] n30759_o;
  wire [23:0] n30760_o;
  wire [23:0] n30761_o;
  wire [23:0] n30762_o;
  wire [23:0] n30763_o;
  wire [23:0] n30764_o;
  wire n30765_o;
  wire n30766_o;
  wire n30767_o;
  wire n30768_o;
  wire n30769_o;
  wire n30770_o;
  wire n30772_o;
  wire [18:0] n30773_o;
  wire n30775_o;
  wire [4:0] n30776_o;
  wire n30778_o;
  wire n30779_o;
  wire [4:0] n30780_o;
  wire [4:0] n30782_o;
  wire n30783_o;
  wire [18:0] n30784_o;
  wire n30786_o;
  wire [4:0] n30787_o;
  wire n30788_o;
  wire n30789_o;
  wire [4:0] n30790_o;
  wire [4:0] n30792_o;
  wire [4:0] n30794_o;
  wire [4:0] n30795_o;
  wire [4:0] n30797_o;
  wire n30798_o;
  wire [4:0] n30801_o;
  wire [4:0] n30802_o;
  wire [4:0] n30805_o;
  wire [2:0] n30828_o;
  wire n30924_o;
  reg [24:0] n31324_burst_min_v;
  wire n31330_o;
  wire n31332_o;
  wire n31333_o;
  wire n31334_o;
  wire n31338_o;
  wire [23:0] n31339_o;
  wire [23:0] n31340_o;
  wire [24:0] n31341_o;
  wire [24:0] n31342_o;
  wire [23:0] n31343_o;
  wire [23:0] n31344_o;
  wire [24:0] n31345_o;
  wire [24:0] n31346_o;
  wire [23:0] n31347_o;
  wire [23:0] n31348_o;
  wire [24:0] n31349_o;
  wire [24:0] n31350_o;
  wire [23:0] n31351_o;
  wire [23:0] n31352_o;
  wire [24:0] n31353_o;
  wire [24:0] n31354_o;
  wire [23:0] n31355_o;
  wire [23:0] n31356_o;
  wire [24:0] n31357_o;
  wire [24:0] n31358_o;
  wire [21:0] n31359_o;
  wire n31360_o;
  wire n31361_o;
  wire n31362_o;
  wire n31363_o;
  wire n31364_o;
  wire n31365_o;
  wire n31366_o;
  wire n31367_o;
  wire n31368_o;
  wire [24:0] n31369_o;
  wire [23:0] n31370_o;
  wire [31:0] n31371_o;
  wire [23:0] n31372_o;
  wire n31374_o;
  wire [20:0] n31375_o;
  wire n31378_o;
  wire [21:0] n31379_o;
  wire n31382_o;
  wire [22:0] n31383_o;
  wire [23:0] n31385_o;
  wire [23:0] n31386_o;
  wire [23:0] n31387_o;
  wire [23:0] n31388_o;
  wire [23:0] n31389_o;
  wire [23:0] n31390_o;
  wire [23:0] n31391_o;
  wire [24:0] n31392_o;
  wire [24:0] n31394_o;
  wire [24:0] n31395_o;
  wire [24:0] n31396_o;
  wire [23:0] n31397_o;
  wire n31399_o;
  wire n31402_o;
  wire n31404_o;
  wire [1:0] n31405_o;
  wire n31407_o;
  wire [1:0] n31408_o;
  wire n31410_o;
  wire [23:0] n31413_o;
  wire [23:0] n31415_o;
  wire n31417_o;
  wire [1:0] n31418_o;
  wire n31420_o;
  wire [1:0] n31421_o;
  wire n31423_o;
  wire [23:0] n31426_o;
  wire [23:0] n31428_o;
  wire n31430_o;
  wire [1:0] n31431_o;
  wire n31433_o;
  wire [1:0] n31434_o;
  wire n31436_o;
  wire [23:0] n31439_o;
  wire [23:0] n31441_o;
  wire [23:0] n31442_o;
  wire [23:0] n31443_o;
  wire [23:0] n31444_o;
  wire [23:0] n31445_o;
  wire [23:0] n31447_o;
  wire [23:0] n31448_o;
  wire [23:0] n31449_o;
  wire [23:0] n31450_o;
  wire [24:0] n31451_o;
  wire [23:0] n31452_o;
  wire [23:0] n31453_o;
  wire [24:0] n31454_o;
  wire [23:0] n31455_o;
  wire [23:0] n31456_o;
  wire [24:0] n31457_o;
  wire [23:0] n31458_o;
  wire [23:0] n31459_o;
  wire [24:0] n31460_o;
  wire [23:0] n31461_o;
  wire [23:0] n31462_o;
  wire [24:0] n31463_o;
  wire [31:0] n31464_o;
  wire [23:0] n31465_o;
  wire [24:0] n31466_o;
  wire [24:0] n31467_o;
  wire [24:0] n31468_o;
  wire [2:0] n31469_o;
  wire [23:0] n31470_o;
  wire n31472_o;
  wire [20:0] n31473_o;
  wire n31476_o;
  wire [21:0] n31477_o;
  wire n31480_o;
  wire [22:0] n31481_o;
  wire [23:0] n31483_o;
  wire [23:0] n31484_o;
  wire [23:0] n31485_o;
  wire [23:0] n31486_o;
  wire [23:0] n31487_o;
  wire [23:0] n31488_o;
  wire [23:0] n31489_o;
  wire [23:0] n31490_o;
  wire n31492_o;
  wire n31495_o;
  wire n31497_o;
  wire [1:0] n31498_o;
  wire n31500_o;
  wire [1:0] n31502_o;
  wire n31504_o;
  wire [23:0] n31507_o;
  wire [23:0] n31508_o;
  wire n31510_o;
  wire [1:0] n31511_o;
  wire n31513_o;
  wire [1:0] n31515_o;
  wire n31517_o;
  wire [23:0] n31520_o;
  wire [23:0] n31521_o;
  wire n31523_o;
  wire [1:0] n31524_o;
  wire n31526_o;
  wire [1:0] n31528_o;
  wire n31530_o;
  wire [23:0] n31533_o;
  wire [23:0] n31534_o;
  wire [23:0] n31535_o;
  wire [23:0] n31536_o;
  wire [23:0] n31537_o;
  wire [23:0] n31538_o;
  wire n31540_o;
  wire n31542_o;
  wire n31544_o;
  wire n31546_o;
  wire n31548_o;
  wire n31549_o;
  wire n31550_o;
  wire n31551_o;
  wire n31552_o;
  wire n31553_o;
  wire n31554_o;
  wire [1:0] n31557_o;
  wire n31558_o;
  wire n31559_o;
  wire n31560_o;
  wire n31561_o;
  wire [1:0] n31564_o;
  wire [1:0] n31566_o;
  wire [1:0] n31567_o;
  wire n31569_o;
  wire [20:0] n31571_o;
  wire [20:0] n31573_o;
  wire n31575_o;
  wire [21:0] n31577_o;
  wire [21:0] n31579_o;
  wire n31581_o;
  wire [22:0] n31583_o;
  wire [22:0] n31585_o;
  wire [23:0] n31587_o;
  wire [23:0] n31588_o;
  wire [23:0] n31589_o;
  wire [23:0] n31590_o;
  wire [23:0] n31591_o;
  wire [23:0] n31592_o;
  wire [23:0] n31593_o;
  wire n31595_o;
  wire n31598_o;
  wire [7:0] n31599_o;
  wire [7:0] n31600_o;
  wire [15:0] n31601_o;
  wire [7:0] n31602_o;
  wire [23:0] n31603_o;
  wire [7:0] n31604_o;
  wire [31:0] n31605_o;
  wire [7:0] n31606_o;
  wire [39:0] n31607_o;
  wire [7:0] n31608_o;
  wire [47:0] n31609_o;
  wire [7:0] n31610_o;
  wire [55:0] n31611_o;
  wire [7:0] n31612_o;
  wire [63:0] n31613_o;
  wire [7:0] n31614_o;
  wire [7:0] n31615_o;
  wire [15:0] n31616_o;
  wire [7:0] n31617_o;
  wire [23:0] n31618_o;
  wire [7:0] n31619_o;
  wire [31:0] n31620_o;
  wire [7:0] n31621_o;
  wire [39:0] n31622_o;
  wire [7:0] n31623_o;
  wire [47:0] n31624_o;
  wire [7:0] n31625_o;
  wire [55:0] n31626_o;
  wire [7:0] n31627_o;
  wire [63:0] n31628_o;
  wire [63:0] n31629_o;
  wire [23:0] n31630_o;
  wire n31632_o;
  wire n31635_o;
  wire [514:0] n31636_o;
  wire [104:0] n31637_o;
  wire [47:0] n31638_o;
  wire [72:0] n31646_o;
  wire [72:0] n31647_o;
  wire [72:0] n31648_o;
  wire [72:0] n31649_o;
  wire [72:0] n31650_o;
  wire [49:0] n31651_o;
  wire [79:0] n31652_o;
  wire [47:0] n31653_o;
  wire [24:0] n31672_o;
  wire [23:0] n31673_o;
  wire n31684_o;
  wire n31685_o;
  wire [24:0] n31703_o;
  wire [24:0] n31706_o;
  wire [24:0] n31707_o;
  wire [24:0] n31708_o;
  wire [24:0] n31709_o;
  wire [24:0] n31710_o;
  wire n31712_o;
  wire n31715_o;
  wire n31716_o;
  wire n31717_o;
  wire [24:0] n31718_o;
  wire n31719_o;
  wire [24:0] n31720_o;
  wire [24:0] n31721_o;
  wire n31722_o;
  wire [24:0] n31723_o;
  wire [24:0] n31724_o;
  wire [24:0] n31725_o;
  wire n31726_o;
  wire [24:0] n31727_o;
  wire [24:0] n31728_o;
  wire [24:0] n31729_o;
  wire [24:0] n31730_o;
  wire n31731_o;
  wire [24:0] n31732_o;
  wire [24:0] n31733_o;
  wire [24:0] n31734_o;
  wire [24:0] n31735_o;
  wire [24:0] n31736_o;
  wire n31737_o;
  wire [24:0] n31738_o;
  wire [24:0] n31739_o;
  wire [24:0] n31740_o;
  wire [24:0] n31741_o;
  wire [24:0] n31742_o;
  wire [24:0] n31743_o;
  wire [23:0] n31745_o;
  wire [23:0] n31747_o;
  wire [24:0] n31748_o;
  wire [24:0] n31749_o;
  wire [24:0] n31750_o;
  wire [24:0] n31751_o;
  wire [24:0] n31752_o;
  wire [24:0] n31753_o;
  wire n31754_o;
  wire [23:0] n31755_o;
  wire [23:0] n31757_o;
  wire [23:0] n31758_o;
  wire [23:0] n31760_o;
  wire [24:0] n31761_o;
  wire [24:0] n31762_o;
  wire [24:0] n31763_o;
  wire [24:0] n31764_o;
  wire [24:0] n31765_o;
  wire [24:0] n31766_o;
  wire n31767_o;
  wire [23:0] n31768_o;
  wire [23:0] n31769_o;
  wire [23:0] n31771_o;
  wire [23:0] n31772_o;
  wire [23:0] n31773_o;
  wire [23:0] n31775_o;
  wire [24:0] n31776_o;
  wire [24:0] n31777_o;
  wire [24:0] n31778_o;
  wire [24:0] n31779_o;
  wire [24:0] n31780_o;
  wire [24:0] n31781_o;
  wire n31782_o;
  wire [23:0] n31783_o;
  wire [23:0] n31784_o;
  wire [23:0] n31785_o;
  wire [23:0] n31787_o;
  wire [23:0] n31788_o;
  wire [23:0] n31789_o;
  wire [23:0] n31790_o;
  wire [23:0] n31792_o;
  wire [24:0] n31793_o;
  wire [24:0] n31794_o;
  wire [24:0] n31795_o;
  wire [24:0] n31796_o;
  wire [24:0] n31797_o;
  wire [24:0] n31798_o;
  wire n31799_o;
  wire [23:0] n31800_o;
  wire [23:0] n31801_o;
  wire [23:0] n31802_o;
  wire [23:0] n31803_o;
  wire [23:0] n31805_o;
  wire [23:0] n31806_o;
  wire [23:0] n31807_o;
  wire [23:0] n31808_o;
  wire [23:0] n31809_o;
  wire [23:0] n31811_o;
  wire [24:0] n31812_o;
  wire [24:0] n31813_o;
  wire [24:0] n31814_o;
  wire [24:0] n31815_o;
  wire [24:0] n31816_o;
  wire [24:0] n31817_o;
  wire n31818_o;
  wire [23:0] n31819_o;
  wire [23:0] n31820_o;
  wire [23:0] n31821_o;
  wire [23:0] n31822_o;
  wire [23:0] n31823_o;
  wire [23:0] n31824_o;
  wire [23:0] n31825_o;
  wire [23:0] n31826_o;
  wire [23:0] n31827_o;
  wire [23:0] n31828_o;
  wire [23:0] n31830_o;
  wire [23:0] n31832_o;
  wire [24:0] n31833_o;
  wire [24:0] n31834_o;
  wire [24:0] n31835_o;
  wire [24:0] n31836_o;
  wire [24:0] n31837_o;
  wire [24:0] n31838_o;
  wire n31839_o;
  wire n31840_o;
  wire n31841_o;
  wire [2:0] n31842_o;
  wire n31844_o;
  wire [23:0] n31845_o;
  wire n31846_o;
  wire n31847_o;
  wire [24:0] n31848_o;
  wire [24:0] n31849_o;
  wire [24:0] n31850_o;
  wire n31851_o;
  wire [2:0] n31853_o;
  wire n31855_o;
  wire [23:0] n31856_o;
  wire n31857_o;
  wire n31858_o;
  wire [24:0] n31859_o;
  wire [24:0] n31860_o;
  wire [24:0] n31861_o;
  wire n31862_o;
  wire [2:0] n31864_o;
  wire n31866_o;
  wire [23:0] n31867_o;
  wire n31868_o;
  wire n31869_o;
  wire [24:0] n31870_o;
  wire [24:0] n31871_o;
  wire [24:0] n31872_o;
  wire n31873_o;
  wire [2:0] n31875_o;
  wire n31877_o;
  wire [23:0] n31878_o;
  wire n31879_o;
  wire n31880_o;
  wire [24:0] n31881_o;
  wire [24:0] n31882_o;
  wire [24:0] n31883_o;
  wire n31884_o;
  wire [2:0] n31886_o;
  wire n31888_o;
  wire [23:0] n31889_o;
  wire n31890_o;
  wire n31891_o;
  wire [24:0] n31892_o;
  wire [24:0] n31893_o;
  wire [24:0] n31894_o;
  wire [23:0] n31897_o;
  wire [23:0] n31899_o;
  wire n31900_o;
  wire [23:0] n31901_o;
  wire [23:0] n31903_o;
  wire [23:0] n31904_o;
  wire [23:0] n31906_o;
  wire [24:0] n31907_o;
  wire [23:0] n31908_o;
  wire [23:0] n31909_o;
  wire [23:0] n31911_o;
  wire [23:0] n31912_o;
  wire [23:0] n31913_o;
  wire [23:0] n31915_o;
  wire [24:0] n31916_o;
  wire [23:0] n31917_o;
  wire [23:0] n31918_o;
  wire [23:0] n31919_o;
  wire [23:0] n31921_o;
  wire [23:0] n31922_o;
  wire [23:0] n31923_o;
  wire [23:0] n31924_o;
  wire [23:0] n31926_o;
  wire [24:0] n31927_o;
  wire [23:0] n31928_o;
  wire [23:0] n31929_o;
  wire [23:0] n31930_o;
  wire [23:0] n31931_o;
  wire [23:0] n31933_o;
  wire [23:0] n31934_o;
  wire [23:0] n31935_o;
  wire [23:0] n31936_o;
  wire [23:0] n31937_o;
  wire [23:0] n31939_o;
  wire [24:0] n31940_o;
  wire [23:0] n31941_o;
  wire [23:0] n31942_o;
  wire [23:0] n31943_o;
  wire [23:0] n31944_o;
  wire [23:0] n31945_o;
  wire [23:0] n31946_o;
  wire [23:0] n31947_o;
  wire [23:0] n31948_o;
  wire [23:0] n31949_o;
  wire [23:0] n31950_o;
  wire [24:0] n31951_o;
  wire [23:0] n31953_o;
  wire [23:0] n31955_o;
  wire n31957_o;
  wire n31959_o;
  wire n31961_o;
  wire [23:0] n31963_o;
  wire [23:0] n31965_o;
  wire [23:0] n31967_o;
  wire [23:0] n31969_o;
  wire [23:0] n31971_o;
  wire [23:0] n31973_o;
  wire [23:0] n31975_o;
  wire [23:0] n31977_o;
  wire [23:0] n31979_o;
  wire [23:0] n31981_o;
  wire [23:0] n31983_o;
  wire [23:0] n31985_o;
  wire [24:0] n31986_o;
  wire [24:0] n31987_o;
  wire [24:0] n31988_o;
  wire [24:0] n31989_o;
  wire [24:0] n31990_o;
  wire n31991_o;
  wire [24:0] n31992_o;
  wire n31994_o;
  wire n31996_o;
  wire n31998_o;
  wire n32000_o;
  wire n32002_o;
  wire n32004_o;
  wire n32006_o;
  wire n32008_o;
  wire n32010_o;
  wire [23:0] n32012_o;
  wire [23:0] n32014_o;
  wire [23:0] n32016_o;
  wire [23:0] n32018_o;
  wire [23:0] n32020_o;
  wire [23:0] n32022_o;
  wire [23:0] n32024_o;
  wire [23:0] n32026_o;
  wire [23:0] n32028_o;
  wire [23:0] n32030_o;
  wire [24:0] n32031_o;
  wire [23:0] n32033_o;
  wire [23:0] n32035_o;
  wire [23:0] n32036_o;
  wire n32039_o;
  wire n32040_o;
  wire n32041_o;
  wire n32042_o;
  wire n32043_o;
  wire n32044_o;
  wire n32045_o;
  wire n32046_o;
  wire n32047_o;
  wire n32048_o;
  wire n32049_o;
  wire n32050_o;
  wire n32051_o;
  wire n32052_o;
  wire n32053_o;
  wire n32054_o;
  wire n32055_o;
  wire n32056_o;
  wire n32057_o;
  wire n32058_o;
  wire n32059_o;
  wire n32060_o;
  wire n32061_o;
  wire n32062_o;
  wire n32063_o;
  wire n32064_o;
  wire n32065_o;
  wire n32066_o;
  wire n32067_o;
  wire n32069_o;
  wire n32074_o;
  wire n32076_o;
  wire n32078_o;
  wire n32096_o;
  wire n32099_o;
  wire n32101_o;
  wire n32103_o;
  wire n32105_o;
  wire n32107_o;
  wire n32109_o;
  wire n32111_o;
  wire n32113_o;
  wire n32115_o;
  wire n32131_o;
  wire n32132_o;
  wire n32133_o;
  wire n32134_o;
  wire n32135_o;
  wire n32136_o;
  wire n32137_o;
  wire n32138_o;
  wire n32139_o;
  wire n32140_o;
  wire n32143_o;
  wire n32144_o;
  wire n32145_o;
  wire n32146_o;
  wire n32147_o;
  wire n32148_o;
  wire n32149_o;
  wire n32150_o;
  wire n32151_o;
  wire n32152_o;
  wire n32153_o;
  wire n32154_o;
  wire n32155_o;
  wire n32156_o;
  wire n32157_o;
  wire n32158_o;
  wire n32159_o;
  wire n32160_o;
  wire n32162_o;
  wire n32164_o;
  wire n32417_o;
  wire n32418_o;
  wire [24:0] n32419_o;
  reg [24:0] n32420_q;
  wire n32429_o;
  wire n32430_o;
  wire [47:0] n32431_o;
  wire [47:0] n32432_o;
  reg [47:0] n32433_q;
  wire n32434_o;
  wire n32435_o;
  wire [104:0] n32436_o;
  wire [104:0] n32437_o;
  reg [104:0] n32438_q;
  wire n32439_o;
  wire n32440_o;
  wire [514:0] n32441_o;
  wire [514:0] n32442_o;
  reg [514:0] n32443_q;
  wire [775:0] n32446_o;
  wire [23:0] n32447_o;
  reg [23:0] n32448_q;
  wire [23:0] n32449_o;
  reg [23:0] n32450_q;
  wire [23:0] n32451_o;
  reg [23:0] n32452_q;
  wire [23:0] n32453_o;
  reg [23:0] n32454_q;
  wire [23:0] n32455_o;
  reg [23:0] n32456_q;
  wire [23:0] n32457_o;
  reg [23:0] n32458_q;
  wire [23:0] n32459_o;
  reg [23:0] n32460_q;
  wire [23:0] n32461_o;
  reg [23:0] n32462_q;
  wire [23:0] n32463_o;
  reg [23:0] n32464_q;
  wire [23:0] n32465_o;
  reg [23:0] n32466_q;
  wire [23:0] n32467_o;
  reg [23:0] n32468_q;
  wire [23:0] n32469_o;
  reg [23:0] n32470_q;
  wire [23:0] n32473_o;
  reg [23:0] n32474_q;
  wire n32475_o;
  reg n32476_q;
  wire [24:0] n32477_o;
  reg [24:0] n32478_q;
  wire [24:0] n32479_o;
  reg [24:0] n32480_q;
  wire [24:0] n32481_o;
  reg [24:0] n32482_q;
  wire [24:0] n32483_o;
  reg [24:0] n32484_q;
  wire [24:0] n32485_o;
  reg [24:0] n32486_q;
  wire [23:0] n32487_o;
  reg [23:0] n32488_q;
  wire [24:0] n32489_o;
  reg [24:0] n32490_q;
  wire [3:0] n32491_o;
  reg [3:0] n32492_q;
  wire [3:0] n32493_o;
  reg [3:0] n32494_q;
  wire [3:0] n32495_o;
  reg [3:0] n32496_q;
  wire [26:0] n32497_o;
  reg [26:0] n32498_q;
  wire [3:0] n32499_o;
  reg [3:0] n32500_q;
  wire [3:0] n32501_o;
  reg [3:0] n32502_q;
  wire [26:0] n32503_o;
  reg [26:0] n32504_q;
  wire [3:0] n32505_o;
  reg [3:0] n32506_q;
  wire [3:0] n32507_o;
  reg [3:0] n32508_q;
  wire n32509_o;
  wire n32510_o;
  wire [47:0] n32511_o;
  wire [47:0] n32512_o;
  reg [47:0] n32513_q;
  wire n32514_o;
  wire n32515_o;
  wire [79:0] n32516_o;
  wire [79:0] n32517_o;
  reg [79:0] n32518_q;
  wire n32519_o;
  wire n32520_o;
  wire [2:0] n32521_o;
  wire [2:0] n32522_o;
  reg [2:0] n32523_q;
  wire n32524_o;
  wire n32525_o;
  wire [49:0] n32526_o;
  wire [49:0] n32527_o;
  reg [49:0] n32528_q;
  wire n32529_o;
  wire n32530_o;
  wire [72:0] n32531_o;
  wire [72:0] n32532_o;
  reg [72:0] n32533_q;
  wire n32534_o;
  wire n32535_o;
  wire [72:0] n32536_o;
  wire [72:0] n32537_o;
  reg [72:0] n32538_q;
  wire n32539_o;
  wire n32540_o;
  wire [72:0] n32541_o;
  wire [72:0] n32542_o;
  reg [72:0] n32543_q;
  wire n32544_o;
  wire n32545_o;
  wire [72:0] n32546_o;
  wire [72:0] n32547_o;
  reg [72:0] n32548_q;
  wire n32549_o;
  wire n32550_o;
  wire [72:0] n32551_o;
  wire [72:0] n32552_o;
  reg [72:0] n32553_q;
  wire [775:0] n32562_o;
  wire [23:0] n32563_o;
  reg [23:0] n32564_q;
  wire [23:0] n32565_o;
  reg [23:0] n32566_q;
  wire [23:0] n32567_o;
  reg [23:0] n32568_q;
  wire [23:0] n32569_o;
  reg [23:0] n32570_q;
  wire [23:0] n32571_o;
  reg [23:0] n32572_q;
  wire [23:0] n32573_o;
  reg [23:0] n32574_q;
  wire [23:0] n32575_o;
  reg [23:0] n32576_q;
  wire [23:0] n32577_o;
  reg [23:0] n32578_q;
  wire [23:0] n32579_o;
  reg [23:0] n32580_q;
  wire [23:0] n32581_o;
  reg [23:0] n32582_q;
  wire [24:0] n32583_o;
  reg [24:0] n32584_q;
  wire [23:0] n32585_o;
  reg [23:0] n32586_q;
  wire [23:0] n32587_o;
  reg [23:0] n32588_q;
  wire [23:0] n32591_o;
  reg [23:0] n32592_q;
  wire n32593_o;
  reg n32594_q;
  wire [23:0] n32595_o;
  reg [23:0] n32596_q;
  wire n32599_o;
  reg n32600_q;
  wire n32601_o;
  reg n32602_q;
  wire n32603_o;
  reg n32604_q;
  wire n32605_o;
  reg n32606_q;
  wire [2:0] n32607_o;
  reg [2:0] n32608_q;
  wire [1:0] n32609_o;
  reg [1:0] n32610_q;
  wire [1:0] n32611_o;
  reg [1:0] n32612_q;
  wire [1:0] n32613_o;
  reg [1:0] n32614_q;
  wire [1:0] n32615_o;
  reg [1:0] n32616_q;
  wire [1:0] n32617_o;
  reg [1:0] n32618_q;
  wire [1:0] n32619_o;
  reg [1:0] n32620_q;
  wire [1:0] n32621_o;
  reg [1:0] n32622_q;
  wire [1:0] n32623_o;
  reg [1:0] n32624_q;
  wire [1:0] n32625_o;
  reg [1:0] n32626_q;
  wire [1:0] n32627_o;
  reg [1:0] n32628_q;
  wire [1:0] n32629_o;
  reg [1:0] n32630_q;
  wire [1:0] n32631_o;
  reg [1:0] n32632_q;
  wire [1:0] n32633_o;
  reg [1:0] n32634_q;
  wire [1:0] n32635_o;
  reg [1:0] n32636_q;
  wire [1:0] n32637_o;
  reg [1:0] n32638_q;
  wire [1:0] n32639_o;
  reg [1:0] n32640_q;
  wire [1:0] n32641_o;
  reg [1:0] n32642_q;
  wire [1:0] n32643_o;
  reg [1:0] n32644_q;
  wire [1:0] n32645_o;
  reg [1:0] n32646_q;
  wire [1:0] n32647_o;
  reg [1:0] n32648_q;
  wire [1:0] n32649_o;
  reg [1:0] n32650_q;
  wire [1:0] n32651_o;
  reg [1:0] n32652_q;
  wire [1:0] n32653_o;
  reg [1:0] n32654_q;
  wire [1:0] n32655_o;
  reg [1:0] n32656_q;
  wire n32657_o;
  reg n32658_q;
  wire n32659_o;
  reg n32660_q;
  wire n32661_o;
  reg n32662_q;
  wire n32663_o;
  reg n32664_q;
  wire [5:0] n32665_o;
  reg [5:0] n32666_q;
  wire [5:0] n32667_o;
  reg [5:0] n32668_q;
  wire [5:0] n32669_o;
  reg [5:0] n32670_q;
  wire [5:0] n32671_o;
  reg [5:0] n32672_q;
  wire [63:0] n32673_o;
  reg [63:0] n32674_q;
  wire [63:0] n32675_o;
  reg [63:0] n32676_q;
  wire [63:0] n32677_o;
  reg [63:0] n32678_q;
  wire [63:0] n32679_o;
  reg [63:0] n32680_q;
  wire [23:0] n32681_o;
  reg [23:0] n32682_q;
  wire [23:0] n32683_o;
  reg [23:0] n32684_q;
  wire [23:0] n32685_o;
  reg [23:0] n32686_q;
  wire [31:0] n32687_o;
  reg [31:0] n32688_q;
  wire [23:0] n32689_o;
  reg [23:0] n32690_q;
  wire [23:0] n32691_o;
  reg [23:0] n32692_q;
  wire [23:0] n32693_o;
  reg [23:0] n32694_q;
  wire [31:0] n32695_o;
  reg [31:0] n32696_q;
  wire [31:0] n32697_o;
  reg [31:0] n32698_q;
  wire [4:0] n32699_o;
  reg [4:0] n32700_q;
  wire [4:0] n32701_o;
  reg [4:0] n32702_q;
  wire n32703_o;
  reg n32704_q;
  wire [23:0] n32705_o;
  reg [23:0] n32706_q;
  wire [23:0] n32707_o;
  reg [23:0] n32708_q;
  wire [23:0] n32709_o;
  reg [23:0] n32710_q;
  wire [31:0] n32711_o;
  reg [31:0] n32712_q;
  wire [23:0] n32713_o;
  reg [23:0] n32714_q;
  wire [23:0] n32715_o;
  reg [23:0] n32716_q;
  wire [23:0] n32717_o;
  reg [23:0] n32718_q;
  wire [31:0] n32719_o;
  reg [31:0] n32720_q;
  wire [31:0] n32721_o;
  reg [31:0] n32722_q;
  wire [4:0] n32723_o;
  reg [4:0] n32724_q;
  wire [4:0] n32725_o;
  reg [4:0] n32726_q;
  wire n32727_o;
  reg n32728_q;
  wire n32729_o;
  reg n32730_q;
  wire n32731_o;
  reg n32732_q;
  wire n32733_o;
  reg n32734_q;
  wire n32735_o;
  reg n32736_q;
  wire n32737_o;
  reg n32738_q;
  wire [1:0] n32739_o;
  reg [1:0] n32740_q;
  wire [1:0] n32741_o;
  reg [1:0] n32742_q;
  wire [1:0] n32743_o;
  reg [1:0] n32744_q;
  wire [1:0] n32745_o;
  reg [1:0] n32746_q;
  wire n32747_o;
  reg n32748_q;
  wire n32749_o;
  reg n32750_q;
  wire n32751_o;
  reg n32752_q;
  wire n32753_o;
  reg n32754_q;
  wire n32755_o;
  reg n32756_q;
  wire n32757_o;
  reg n32758_q;
  wire n32759_o;
  reg n32760_q;
  wire n32761_o;
  reg n32762_q;
  wire n32763_o;
  reg n32764_q;
  wire n32765_o;
  reg n32766_q;
  wire n32767_o;
  reg n32768_q;
  wire n32769_o;
  reg n32770_q;
  wire [1:0] n32771_o;
  reg [1:0] n32772_q;
  wire [1:0] n32773_o;
  reg [1:0] n32774_q;
  wire [1:0] n32775_o;
  reg [1:0] n32776_q;
  wire [1:0] n32777_o;
  reg [1:0] n32778_q;
  wire n32779_o;
  reg n32780_q;
  wire n32781_o;
  reg n32782_q;
  wire n32783_o;
  reg n32784_q;
  wire n32787_o;
  reg n32788_q;
  wire n32789_o;
  reg n32790_q;
  wire n32791_o;
  reg n32792_q;
  wire [2:0] n32795_o;
  reg [2:0] n32796_q;
  wire [2:0] n32797_o;
  reg [2:0] n32798_q;
  wire [2:0] n32799_o;
  reg [2:0] n32800_q;
  wire [2:0] n32801_o;
  reg [2:0] n32802_q;
  wire [2:0] n32803_o;
  reg [2:0] n32804_q;
  wire [2:0] n32805_o;
  reg [2:0] n32806_q;
  wire [2:0] n32807_o;
  reg [2:0] n32808_q;
  wire [2:0] n32809_o;
  reg [2:0] n32810_q;
  wire n32811_o;
  reg n32812_q;
  wire n32813_o;
  reg n32814_q;
  wire n32815_o;
  reg n32816_q;
  wire n32817_o;
  reg n32818_q;
  wire n32819_o;
  reg n32820_q;
  wire n32821_o;
  reg n32822_q;
  wire n32823_o;
  reg n32824_q;
  wire n32825_o;
  reg n32826_q;
  wire [1:0] n32827_o;
  reg [1:0] n32828_q;
  wire [1:0] n32829_o;
  reg [1:0] n32830_q;
  wire [1:0] n32831_o;
  reg [1:0] n32832_q;
  wire [1:0] n32833_o;
  reg [1:0] n32834_q;
  wire [1:0] n32835_o;
  reg [1:0] n32836_q;
  wire [1:0] n32837_o;
  reg [1:0] n32838_q;
  wire [1:0] n32839_o;
  reg [1:0] n32840_q;
  wire [1:0] n32841_o;
  reg [1:0] n32842_q;
  wire n32843_o;
  reg n32844_q;
  wire n32845_o;
  reg n32846_q;
  wire n32847_o;
  reg n32848_q;
  wire n32849_o;
  reg n32850_q;
  reg [2:0] n32852_q;
  reg [2:0] n32853_q;
  reg [5:0] n32854_q;
  reg [5:0] n32855_q;
  wire [24:0] n32856_o;
  reg [24:0] n32857_q;
  wire [31:0] n32858_o;
  wire [31:0] n32859_o;
  reg [31:0] n32860_q;
  reg n32861_q;
  reg n32864_q;
  wire n32865_o;
  wire n32866_o;
  wire n32867_o;
  wire n32868_o;
  wire n32869_o;
  wire n32870_o;
  wire n32871_o;
  wire [4:0] n32872_o;
  wire [4:0] n32873_o;
  wire [4:0] n32874_o;
  wire n32875_o;
  wire [4:0] n32876_o;
  wire n32877_o;
  wire [4:0] n32878_o;
  wire [4:0] n32879_o;
  wire [4:0] n32880_o;
  wire [4:0] n32881_o;
  wire n32882_o;
  wire [4:0] n32883_o;
  wire n32884_o;
  wire [4:0] n32885_o;
  wire n32886_o;
  wire n32887_o;
  wire n32888_o;
  wire n32889_o;
  wire n32890_o;
  wire n32891_o;
  wire n32892_o;
  assign ready_out = ready;
  assign gen_valid_out = gen_valid_r;
  assign gen_vm_out = vm_rrrr;
  assign gen_fork_out = n30331_o;
  assign gen_data_flow_out = data_flow_rrrr;
  assign gen_src_stream_out = stream_src_rrrr;
  assign gen_dest_stream_out = stream_dest_rrrr;
  assign gen_stream_id_out = stream_id_rrrr;
  assign gen_src_vector_out = src_vector_rrrr;
  assign gen_dst_vector_out = dst_vector_rrrr;
  assign gen_src_scatter_out = src_scatter_rrrr;
  assign gen_dst_scatter_out = dst_scatter_rrrr;
  assign gen_src_start_out = s_burstpos_start_rrrr;
  assign gen_src_end_out = s_burstpos_end_rrr;
  assign gen_dst_end_out = d_burstpos_end_rrr;
  assign gen_addr_source_out = s_gen_addr_r;
  assign gen_addr_source_mode_out = src_addr_mode_rrrr;
  assign gen_addr_dest_out = d_gen_addr_r;
  assign gen_addr_dest_mode_out = dst_addr_mode_rrrr;
  assign gen_eof_out = n30335_o;
  assign gen_bus_id_source_out = dp_src_bus_id_rrrr;
  assign gen_data_type_source_out = dp_src_data_type_rrrr;
  assign gen_data_model_source_out = dp_src_data_model_rrrr;
  assign gen_bus_id_dest_out = dp_dst_bus_id_rrrr;
  assign gen_busy_dest_out = gen_busy_dest_r;
  assign gen_data_type_dest_out = dp_dst_data_type_rrrr;
  assign gen_data_model_dest_out = dp_dst_data_model_rrrr;
  assign gen_burstlen_source_out = s_gen_burstlen_rr;
  assign gen_burstlen_dest_out = d_gen_burstlen_rr;
  assign gen_thread_out = dp_thread_rrrr;
  assign gen_mcast_out = dp_mcast_rrrr;
  assign gen_data_out = data_rrrr;
  assign log_out = log_r;
  assign log_valid_out = log_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:96:16  */
  assign n29602_o = {instruction_source_in_burst_max_len, instruction_source_in_bufsize, instruction_source_in_bus_id, instruction_source_in_datatype, instruction_source_in_repeat, instruction_source_in_data, instruction_source_in_mcast, instruction_source_in_totalcount, instruction_source_in_scatter, instruction_source_in_data_model, instruction_source_in_double_precision, instruction_source_in_burststride, instruction_source_in_count, instruction_source_in_bar, instruction_source_in_burst_min, instruction_source_in_burst_max_index, instruction_source_in_burst_max_init, instruction_source_in_burst_max2, instruction_source_in_burst_max, instruction_source_in_stride4_min, instruction_source_in_stride4_max, instruction_source_in_stride4_count, instruction_source_in_stride4, instruction_source_in_stride3_min, instruction_source_in_stride3_max, instruction_source_in_stride3_count, instruction_source_in_stride3, instruction_source_in_stride2_min, instruction_source_in_stride2_max, instruction_source_in_stride2_count, instruction_source_in_stride2, instruction_source_in_stride1_min, instruction_source_in_stride1_max, instruction_source_in_stride1_count, instruction_source_in_stride1, instruction_source_in_stride0_min, instruction_source_in_stride0_max, instruction_source_in_stride0_count, instruction_source_in_stride0};
  /* ../../HW/src/dp/dp_gen.vhd:95:16  */
  assign n29603_o = {instruction_dest_in_burst_max_len, instruction_dest_in_bufsize, instruction_dest_in_bus_id, instruction_dest_in_datatype, instruction_dest_in_repeat, instruction_dest_in_data, instruction_dest_in_mcast, instruction_dest_in_totalcount, instruction_dest_in_scatter, instruction_dest_in_data_model, instruction_dest_in_double_precision, instruction_dest_in_burststride, instruction_dest_in_count, instruction_dest_in_bar, instruction_dest_in_burst_min, instruction_dest_in_burst_max_index, instruction_dest_in_burst_max_init, instruction_dest_in_burst_max2, instruction_dest_in_burst_max, instruction_dest_in_stride4_min, instruction_dest_in_stride4_max, instruction_dest_in_stride4_count, instruction_dest_in_stride4, instruction_dest_in_stride3_min, instruction_dest_in_stride3_max, instruction_dest_in_stride3_count, instruction_dest_in_stride3, instruction_dest_in_stride2_min, instruction_dest_in_stride2_max, instruction_dest_in_stride2_count, instruction_dest_in_stride2, instruction_dest_in_stride1_min, instruction_dest_in_stride1_max, instruction_dest_in_stride1_count, instruction_dest_in_stride1, instruction_dest_in_stride0_min, instruction_dest_in_stride0_max, instruction_dest_in_stride0_count, instruction_dest_in_stride0};
  /* ../../HW/src/dp/dp_gen.vhd:94:16  */
  assign n29604_o = {pre_instruction_source_in_burst_max_len, pre_instruction_source_in_bufsize, pre_instruction_source_in_bus_id, pre_instruction_source_in_datatype, pre_instruction_source_in_repeat, pre_instruction_source_in_data, pre_instruction_source_in_mcast, pre_instruction_source_in_totalcount, pre_instruction_source_in_scatter, pre_instruction_source_in_data_model, pre_instruction_source_in_double_precision, pre_instruction_source_in_burststride, pre_instruction_source_in_count, pre_instruction_source_in_bar, pre_instruction_source_in_burst_min, pre_instruction_source_in_burst_max_index, pre_instruction_source_in_burst_max_init, pre_instruction_source_in_burst_max2, pre_instruction_source_in_burst_max, pre_instruction_source_in_stride4_min, pre_instruction_source_in_stride4_max, pre_instruction_source_in_stride4_count, pre_instruction_source_in_stride4, pre_instruction_source_in_stride3_min, pre_instruction_source_in_stride3_max, pre_instruction_source_in_stride3_count, pre_instruction_source_in_stride3, pre_instruction_source_in_stride2_min, pre_instruction_source_in_stride2_max, pre_instruction_source_in_stride2_count, pre_instruction_source_in_stride2, pre_instruction_source_in_stride1_min, pre_instruction_source_in_stride1_max, pre_instruction_source_in_stride1_count, pre_instruction_source_in_stride1, pre_instruction_source_in_stride0_min, pre_instruction_source_in_stride0_max, pre_instruction_source_in_stride0_count, pre_instruction_source_in_stride0};
  /* ../../HW/src/dp/dp_gen.vhd:93:16  */
  assign n29605_o = {pre_instruction_dest_in_burst_max_len, pre_instruction_dest_in_bufsize, pre_instruction_dest_in_bus_id, pre_instruction_dest_in_datatype, pre_instruction_dest_in_repeat, pre_instruction_dest_in_data, pre_instruction_dest_in_mcast, pre_instruction_dest_in_totalcount, pre_instruction_dest_in_scatter, pre_instruction_dest_in_data_model, pre_instruction_dest_in_double_precision, pre_instruction_dest_in_burststride, pre_instruction_dest_in_count, pre_instruction_dest_in_bar, pre_instruction_dest_in_burst_min, pre_instruction_dest_in_burst_max_index, pre_instruction_dest_in_burst_max_init, pre_instruction_dest_in_burst_max2, pre_instruction_dest_in_burst_max, pre_instruction_dest_in_stride4_min, pre_instruction_dest_in_stride4_max, pre_instruction_dest_in_stride4_count, pre_instruction_dest_in_stride4, pre_instruction_dest_in_stride3_min, pre_instruction_dest_in_stride3_max, pre_instruction_dest_in_stride3_count, pre_instruction_dest_in_stride3, pre_instruction_dest_in_stride2_min, pre_instruction_dest_in_stride2_max, pre_instruction_dest_in_stride2_count, pre_instruction_dest_in_stride2, pre_instruction_dest_in_stride1_min, pre_instruction_dest_in_stride1_max, pre_instruction_dest_in_stride1_count, pre_instruction_dest_in_stride1, pre_instruction_dest_in_stride0_min, pre_instruction_dest_in_stride0_max, pre_instruction_dest_in_stride0_count, pre_instruction_dest_in_stride0};
  /* ../../HW/src/dp/dp_gen.vhd:130:8  */
  assign s_template_r = n32446_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:131:8  */
  assign s_i0_r = n32448_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:132:8  */
  assign s_i1_r = n32450_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:133:8  */
  assign s_i2_r = n32452_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:134:8  */
  assign s_i3_r = n32454_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:135:8  */
  assign s_i4_r = n32456_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:136:8  */
  assign s_i0_count_r = n32458_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:137:8  */
  assign s_i1_count_r = n32460_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:138:8  */
  assign s_i2_count_r = n32462_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:139:8  */
  assign s_i3_count_r = n32464_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:140:8  */
  assign s_i4_count_r = n32466_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:141:8  */
  assign s_burstlen_r = n32468_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:142:8  */
  assign s_burstpos_r = n32470_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:144:8  */
  always @*
    s_burstremain_r = n32474_q; // (isignal)
  initial
    s_burstremain_r = 24'b111111111111111111111111;
  /* ../../HW/src/dp/dp_gen.vhd:145:8  */
  always @*
    s_valid_r = n32476_q; // (isignal)
  initial
    s_valid_r = 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:147:8  */
  assign s_i0_start_r = n32478_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:148:8  */
  assign s_i1_start_r = n32480_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:149:8  */
  assign s_i2_start_r = n32482_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:150:8  */
  assign s_i3_start_r = n32484_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:151:8  */
  assign s_i4_start_r = n32486_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:153:8  */
  assign s_burstpos_stride_r = n32488_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:154:8  */
  assign s_burstpos_start_r = n32490_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:155:8  */
  assign s_burstpos_start_rr = n32492_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:156:8  */
  assign s_burstpos_start_rrr = n32494_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:157:8  */
  assign s_burstpos_start_rrrr = n32496_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:159:8  */
  assign s_burstpos_end_r = n32498_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:160:8  */
  assign s_burstpos_end_rr = n32500_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:161:8  */
  assign s_burstpos_end_rrr = n32502_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:163:8  */
  assign d_burstpos_end_r = n32504_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:164:8  */
  assign d_burstpos_end_rr = n32506_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:165:8  */
  assign d_burstpos_end_rrr = n32508_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:168:8  */
  assign d_template_r = n32562_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:169:8  */
  assign d_i0_r = n32564_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:170:8  */
  assign d_i1_r = n32566_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:171:8  */
  assign d_i2_r = n32568_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:172:8  */
  assign d_i3_r = n32570_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:173:8  */
  assign d_i4_r = n32572_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:174:8  */
  assign d_i0_count_r = n32574_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:175:8  */
  assign d_i1_count_r = n32576_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:176:8  */
  assign d_i2_count_r = n32578_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:177:8  */
  assign d_i3_count_r = n32580_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:178:8  */
  assign d_i4_count_r = n32582_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:179:8  */
  assign d_burst_max_r = n32584_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:180:8  */
  assign d_burstlen_r = n32586_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:181:8  */
  assign d_burstpos_r = n32588_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:183:8  */
  always @*
    d_burstremain_r = n32592_q; // (isignal)
  initial
    d_burstremain_r = 24'b111111111111111111111111;
  /* ../../HW/src/dp/dp_gen.vhd:184:8  */
  always @*
    d_valid_r = n32594_q; // (isignal)
  initial
    d_valid_r = 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:186:8  */
  assign currlen_r = n32596_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:187:8  */
  assign currlen_new = n29675_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:189:8  */
  assign reload = n29672_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:191:8  */
  assign s_burstlen_wrap = n30346_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:192:8  */
  assign s_i0_wrap = n30351_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:193:8  */
  assign s_i1_wrap = n30356_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:194:8  */
  assign s_i2_wrap = n30361_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:195:8  */
  assign s_i3_wrap = n30366_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:196:8  */
  assign s_i4_wrap = n30371_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:197:8  */
  assign s_burstlen_new = n30241_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:198:8  */
  assign s_burstpos_new = n30243_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:199:8  */
  assign s_i0_new = n30245_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:200:8  */
  assign s_i1_new = n30247_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:201:8  */
  assign s_i2_new = n30249_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:202:8  */
  assign s_i3_new = n30251_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:203:8  */
  assign s_i4_new = n30253_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:204:8  */
  assign s_i0_count_new = n30278_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:205:8  */
  assign s_i1_count_new = n30280_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:206:8  */
  assign s_i2_count_new = n30282_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:207:8  */
  assign s_i3_count_new = n30284_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:208:8  */
  assign s_i4_count_new = n30286_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:210:8  */
  assign s_burstpos_start_new = n30256_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:211:8  */
  assign s_i0_start_new = n30260_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:212:8  */
  assign s_i1_start_new = n30264_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:213:8  */
  assign s_i2_start_new = n30268_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:214:8  */
  assign s_i3_start_new = n30272_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:215:8  */
  assign s_i4_start_new = n30276_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:217:8  */
  assign d_burstlen_wrap = n30441_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:218:8  */
  assign d_i0_wrap = n30446_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:219:8  */
  assign d_i1_wrap = n30451_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:220:8  */
  assign d_i2_wrap = n30456_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:221:8  */
  assign d_i3_wrap = n30461_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:222:8  */
  assign d_i4_wrap = n30466_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:223:8  */
  assign d_burstlen_new = n30288_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:224:8  */
  assign d_burstpos_new = n30290_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:225:8  */
  assign d_i0_new = n30292_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:226:8  */
  assign d_i1_new = n30294_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:227:8  */
  assign d_i2_new = n30296_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:228:8  */
  assign d_i3_new = n30298_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:229:8  */
  assign d_i4_new = n30300_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:230:8  */
  assign d_i0_new2 = n30304_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:231:8  */
  assign d_i1_new2 = n30308_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:232:8  */
  assign d_i2_new2 = n30312_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:233:8  */
  assign d_i3_new2 = n30316_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:234:8  */
  assign d_i4_new2 = n30320_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:235:8  */
  assign d_i0_count_new = n30322_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:236:8  */
  assign d_i1_count_new = n30324_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:237:8  */
  assign d_i2_count_new = n30326_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:238:8  */
  assign d_i3_count_new = n30328_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:239:8  */
  assign d_i4_count_new = n30330_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:241:8  */
  assign running_r = n32600_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:242:8  */
  assign running_rr = n32602_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:243:8  */
  assign running_rrr = n32604_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:244:8  */
  assign running_rrrr = n32606_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:245:8  */
  assign gen_valid_r = n32608_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:246:8  */
  assign dp_dst_bus_id_r = n32610_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:247:8  */
  assign dp_dst_bus_id_rr = n32612_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:248:8  */
  assign dp_dst_bus_id_rrr = n32614_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:249:8  */
  assign dp_dst_bus_id_rrrr = n32616_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:250:8  */
  assign dp_src_bus_id_r = n32618_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:251:8  */
  assign dp_src_bus_id_rr = n32620_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:252:8  */
  assign dp_src_bus_id_rrr = n32622_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:253:8  */
  assign dp_src_bus_id_rrrr = n32624_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:254:8  */
  assign dp_dst_data_type_r = n32626_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:255:8  */
  assign dp_dst_data_type_rr = n32628_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:256:8  */
  assign dp_dst_data_type_rrr = n32630_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:257:8  */
  assign dp_dst_data_type_rrrr = n32632_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:258:8  */
  assign dp_src_data_type_r = n32634_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:259:8  */
  assign dp_src_data_type_rr = n32636_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:260:8  */
  assign dp_src_data_type_rrr = n32638_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:261:8  */
  assign dp_src_data_type_rrrr = n32640_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:262:8  */
  assign dp_src_data_model_r = n32642_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:263:8  */
  assign dp_src_data_model_rr = n32644_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:264:8  */
  assign dp_src_data_model_rrr = n32646_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:265:8  */
  assign dp_src_data_model_rrrr = n32648_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:266:8  */
  assign dp_dst_data_model_r = n32650_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:267:8  */
  assign dp_dst_data_model_rr = n32652_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:268:8  */
  assign dp_dst_data_model_rrr = n32654_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:269:8  */
  assign dp_dst_data_model_rrrr = n32656_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:270:8  */
  assign dp_thread_r = n32658_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:271:8  */
  assign dp_thread_rr = n32660_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:272:8  */
  assign dp_thread_rrr = n32662_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:273:8  */
  assign dp_thread_rrrr = n32664_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:274:8  */
  always @*
    dp_mcast_r = n32666_q; // (isignal)
  initial
    dp_mcast_r = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:275:8  */
  always @*
    dp_mcast_rr = n32668_q; // (isignal)
  initial
    dp_mcast_rr = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:276:8  */
  always @*
    dp_mcast_rrr = n32670_q; // (isignal)
  initial
    dp_mcast_rrr = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:277:8  */
  always @*
    dp_mcast_rrrr = n32672_q; // (isignal)
  initial
    dp_mcast_rrrr = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:278:8  */
  assign data_r = n32674_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:279:8  */
  assign data_rr = n32676_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:280:8  */
  assign data_rrr = n32678_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:281:8  */
  assign data_rrrr = n32680_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:283:8  */
  assign s_bufsize_r = n32682_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:284:8  */
  assign s_bufsize_rr = n32684_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:285:8  */
  assign s_temp1_r = n32686_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:286:8  */
  assign s_temp2_r = n32688_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:287:8  */
  assign s_temp3_r = n32690_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:288:8  */
  assign s_temp4_r = n32692_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:289:8  */
  assign s_temp5_r = n32694_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:290:8  */
  assign s_temp4_rr = n32696_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:291:8  */
  assign s_gen_addr_r = n32698_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:292:8  */
  assign s_gen_burstlen_r = n32700_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:293:8  */
  assign s_gen_burstlen_rr = n32702_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:294:8  */
  assign s_gen_burstlen_progress_r = n32704_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:296:8  */
  assign s_i0_valid = n30379_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:297:8  */
  assign s_i1_valid = n30387_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:298:8  */
  assign s_i2_valid = n30395_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:299:8  */
  assign s_i3_valid = n30403_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:300:8  */
  assign s_i4_valid = n30411_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:301:8  */
  assign s_burst_valid = n30419_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:303:8  */
  assign s_i0_start_valid = n30422_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:304:8  */
  assign s_i1_start_valid = n30424_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:305:8  */
  assign s_i2_start_valid = n30426_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:306:8  */
  assign s_i3_start_valid = n30428_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:307:8  */
  assign s_i4_start_valid = n30430_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:308:8  */
  assign s_burst_start_valid = n30436_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:310:8  */
  assign d_bufsize_r = n32706_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:311:8  */
  assign d_bufsize_rr = n32708_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:312:8  */
  assign d_temp1_r = n32710_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:313:8  */
  assign d_temp2_r = n32712_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:314:8  */
  assign d_temp3_r = n32714_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:315:8  */
  assign d_temp4_r = n32716_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:316:8  */
  assign d_temp5_r = n32718_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:317:8  */
  assign d_temp4_rr = n32720_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:318:8  */
  assign d_gen_addr_r = n32722_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:319:8  */
  assign d_gen_burstlen_r = n32724_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:320:8  */
  assign d_gen_burstlen_rr = n32726_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:322:8  */
  assign d_i0_valid = n30474_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:323:8  */
  assign d_i1_valid = n30482_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:324:8  */
  assign d_i2_valid = n30490_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:325:8  */
  assign d_i3_valid = n30498_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:326:8  */
  assign d_i4_valid = n30506_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:327:8  */
  assign d_burst_valid = n30514_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:329:8  */
  assign eof_r = n32728_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:330:8  */
  assign eof_rr = n32730_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:331:8  */
  assign eof_rrr = n32732_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:332:8  */
  assign eof_rrrr = n32734_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:333:8  */
  always @*
    done_r = n32736_q; // (isignal)
  initial
    done_r = 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:335:8  */
  assign repeat_r = n32738_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:337:8  */
  assign data_flow_r = n32740_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:338:8  */
  assign data_flow_rr = n32742_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:339:8  */
  assign data_flow_rrr = n32744_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:340:8  */
  assign data_flow_rrrr = n32746_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:342:8  */
  assign stream_src_r = n32748_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:343:8  */
  assign stream_src_rr = n32750_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:344:8  */
  assign stream_src_rrr = n32752_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:345:8  */
  assign stream_src_rrrr = n32754_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:347:8  */
  assign stream_dest_r = n32756_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:348:8  */
  assign stream_dest_rr = n32758_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:349:8  */
  assign stream_dest_rrr = n32760_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:350:8  */
  assign stream_dest_rrrr = n32762_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:352:8  */
  assign vm_r = n32764_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:353:8  */
  assign vm_rr = n32766_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:354:8  */
  assign vm_rrr = n32768_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:355:8  */
  assign vm_rrrr = n32770_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:357:8  */
  assign stream_id_r = n32772_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:358:8  */
  assign stream_id_rr = n32774_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:359:8  */
  assign stream_id_rrr = n32776_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:360:8  */
  assign stream_id_rrrr = n32778_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:362:8  */
  assign src_double_r = n32780_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:363:8  */
  assign src_double_rr = n32782_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:364:8  */
  assign src_double_rrr = n32784_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:367:8  */
  assign dst_double_r = n32788_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:368:8  */
  assign dst_double_rr = n32790_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:369:8  */
  assign dst_double_rrr = n32792_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:372:8  */
  assign src_vector_r = n32796_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:373:8  */
  assign src_vector_rr = n32798_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:374:8  */
  assign src_vector_rrr = n32800_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:375:8  */
  assign src_vector_rrrr = n32802_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:377:8  */
  assign dst_vector_r = n32804_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:378:8  */
  assign dst_vector_rr = n32806_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:379:8  */
  assign dst_vector_rrr = n32808_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:380:8  */
  assign dst_vector_rrrr = n32810_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:382:8  */
  assign src_addr_mode_r = n32812_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:383:8  */
  assign src_addr_mode_rr = n32814_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:384:8  */
  assign src_addr_mode_rrr = n32816_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:385:8  */
  assign src_addr_mode_rrrr = n32818_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:387:8  */
  assign dst_addr_mode_r = n32820_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:388:8  */
  assign dst_addr_mode_rr = n32822_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:389:8  */
  assign dst_addr_mode_rrr = n32824_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:390:8  */
  assign dst_addr_mode_rrrr = n32826_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:392:8  */
  assign src_scatter_r = n32828_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:393:8  */
  assign src_scatter_rr = n32830_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:394:8  */
  assign src_scatter_rrr = n32832_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:395:8  */
  assign src_scatter_rrrr = n32834_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:397:8  */
  assign dst_scatter_r = n32836_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:398:8  */
  assign dst_scatter_rr = n32838_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:399:8  */
  assign dst_scatter_rrr = n32840_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:400:8  */
  assign dst_scatter_rrrr = n32842_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:402:8  */
  assign src_vector = n30234_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:403:8  */
  assign dst_vector = n30236_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:404:8  */
  assign src_scatter = n30237_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:405:8  */
  assign dst_scatter = n30238_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:407:8  */
  assign src_is_burst_r = n32844_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:408:8  */
  assign src_is_burst_rr = n32846_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:409:8  */
  assign dst_is_burst_r = n32848_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:410:8  */
  assign dst_is_burst_rr = n32850_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:413:8  */
  assign src_is_vector_r = n32852_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:414:8  */
  assign dst_is_vector_r = n32853_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:415:8  */
  assign src_is_scatter_r = n32854_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:416:8  */
  assign dst_is_scatter_r = n32855_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:418:8  */
  assign s_burst_actual_max_r = n32857_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:420:8  */
  assign log = n32858_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:421:8  */
  assign log_r = n32860_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:422:8  */
  assign log_valid_r = n32861_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:424:8  */
  assign source_double_precision = n29651_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:425:8  */
  assign dest_double_precision = n29656_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:427:8  */
  assign waitreq = n30341_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:429:8  */
  assign ready = n29667_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:441:8  */
  assign gen_busy_dest_r = n32864_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:452:50  */
  assign n29648_o = n29602_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:452:100  */
  assign n29650_o = instruction_bus_id_source_in != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:452:67  */
  assign n29651_o = n29650_o ? n29648_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:453:46  */
  assign n29653_o = n29603_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:453:94  */
  assign n29655_o = instruction_bus_id_dest_in != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:453:63  */
  assign n29656_o = n29655_o ? n29653_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:456:29  */
  assign n29659_o = ~running_r;
  /* ../../HW/src/dp/dp_gen.vhd:456:48  */
  assign n29660_o = ~running_rr;
  /* ../../HW/src/dp/dp_gen.vhd:456:34  */
  assign n29661_o = n29660_o & n29659_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:68  */
  assign n29662_o = ~running_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:456:53  */
  assign n29663_o = n29662_o & n29661_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:89  */
  assign n29664_o = ~running_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:456:73  */
  assign n29665_o = n29664_o & n29663_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:95  */
  assign n29666_o = reload & n29665_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:14  */
  assign n29667_o = n29666_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:459:30  */
  assign n29670_o = ~running_r;
  /* ../../HW/src/dp/dp_gen.vhd:459:35  */
  assign n29671_o = n29670_o | done_r;
  /* ../../HW/src/dp/dp_gen.vhd:459:15  */
  assign n29672_o = n29671_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:462:25  */
  assign n29675_o = currlen_r - 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:531:12  */
  assign n29686_o = ~reset_in;
  /* ../../HW/src/dp/dp_gen.vhd:541:42  */
  assign n29688_o = n29604_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:541:62  */
  assign n29690_o = n29688_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:542:43  */
  assign n29692_o = pre_instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:541:98  */
  assign n29693_o = n29692_o & n29690_o;
  /* ../../HW/src/dp/dp_gen.vhd:543:37  */
  assign n29694_o = n29604_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:542:98  */
  assign n29695_o = n29694_o & n29693_o;
  /* ../../HW/src/dp/dp_gen.vhd:544:39  */
  assign n29696_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:544:50  */
  assign n29698_o = n29696_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:546:42  */
  assign n29700_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:546:53  */
  assign n29702_o = n29700_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:546:10  */
  assign n29705_o = n29702_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:544:10  */
  assign n29706_o = n29698_o ? 2'b01 : n29705_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:7  */
  assign n29707_o = n29695_o ? n29706_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:40  */
  assign n29708_o = n29605_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:555:60  */
  assign n29710_o = n29708_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:556:41  */
  assign n29712_o = pre_instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:96  */
  assign n29713_o = n29712_o & n29710_o;
  /* ../../HW/src/dp/dp_gen.vhd:557:35  */
  assign n29714_o = n29605_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:556:96  */
  assign n29715_o = n29714_o & n29713_o;
  /* ../../HW/src/dp/dp_gen.vhd:558:37  */
  assign n29716_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:558:48  */
  assign n29718_o = n29716_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:560:40  */
  assign n29719_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:560:51  */
  assign n29721_o = n29719_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:560:10  */
  assign n29722_o = n29721_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:558:10  */
  assign n29723_o = n29718_o ? 2'b01 : n29722_o;
  /* ../../HW/src/dp/dp_gen.vhd:555:7  */
  assign n29724_o = n29715_o ? n29723_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:569:42  */
  assign n29726_o = pre_instruction_bus_id_source_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:570:39  */
  assign n29727_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:570:50  */
  assign n29729_o = n29727_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:571:39  */
  assign n29730_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:571:50  */
  assign n29732_o = n29730_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:572:44  */
  assign n29733_o = n29604_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:572:64  */
  assign n29735_o = n29733_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:571:111  */
  assign n29736_o = n29735_o & n29732_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:111  */
  assign n29737_o = n29729_o | n29736_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:10  */
  assign n29740_o = n29737_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:577:39  */
  assign n29741_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:577:50  */
  assign n29743_o = n29741_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:578:46  */
  assign n29744_o = n29604_o[2:0];
  /* ../../HW/src/dp/dp_gen.vhd:578:66  */
  assign n29746_o = n29744_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:579:46  */
  assign n29747_o = n29604_o[100:98];
  /* ../../HW/src/dp/dp_gen.vhd:579:66  */
  assign n29749_o = n29747_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:578:90  */
  assign n29750_o = n29749_o & n29746_o;
  /* ../../HW/src/dp/dp_gen.vhd:580:46  */
  assign n29751_o = n29604_o[198:196];
  /* ../../HW/src/dp/dp_gen.vhd:580:66  */
  assign n29753_o = n29751_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:579:90  */
  assign n29754_o = n29753_o & n29750_o;
  /* ../../HW/src/dp/dp_gen.vhd:581:46  */
  assign n29755_o = n29604_o[296:294];
  /* ../../HW/src/dp/dp_gen.vhd:581:66  */
  assign n29757_o = n29755_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:580:90  */
  assign n29758_o = n29757_o & n29754_o;
  /* ../../HW/src/dp/dp_gen.vhd:582:46  */
  assign n29759_o = n29604_o[394:392];
  /* ../../HW/src/dp/dp_gen.vhd:582:66  */
  assign n29761_o = n29759_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:581:90  */
  assign n29762_o = n29761_o & n29758_o;
  /* ../../HW/src/dp/dp_gen.vhd:583:39  */
  assign n29763_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:583:50  */
  assign n29765_o = n29763_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:582:90  */
  assign n29766_o = n29765_o & n29762_o;
  /* ../../HW/src/dp/dp_gen.vhd:584:44  */
  assign n29767_o = n29604_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:584:64  */
  assign n29769_o = n29767_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:583:111  */
  assign n29770_o = n29769_o & n29766_o;
  /* ../../HW/src/dp/dp_gen.vhd:585:48  */
  assign n29771_o = n29604_o[492:490];
  /* ../../HW/src/dp/dp_gen.vhd:585:68  */
  assign n29773_o = n29771_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:584:99  */
  assign n29774_o = n29773_o & n29770_o;
  /* ../../HW/src/dp/dp_gen.vhd:586:42  */
  assign n29775_o = n29604_o[595:593];
  /* ../../HW/src/dp/dp_gen.vhd:586:62  */
  assign n29777_o = n29775_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:585:103  */
  assign n29778_o = n29777_o & n29774_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:111  */
  assign n29779_o = n29743_o | n29778_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:7  */
  assign n29782_o = n29779_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:569:7  */
  assign n29783_o = n29726_o ? n29740_o : n29782_o;
  /* ../../HW/src/dp/dp_gen.vhd:593:41  */
  assign n29785_o = pre_instruction_bus_id_dest_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:594:38  */
  assign n29786_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:594:49  */
  assign n29788_o = n29786_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:595:38  */
  assign n29789_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:595:49  */
  assign n29791_o = n29789_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:596:43  */
  assign n29792_o = n29605_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:596:63  */
  assign n29794_o = n29792_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:595:108  */
  assign n29795_o = n29794_o & n29791_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:108  */
  assign n29796_o = n29788_o | n29795_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:11  */
  assign n29799_o = n29796_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:601:35  */
  assign n29800_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:601:46  */
  assign n29802_o = n29800_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:602:42  */
  assign n29803_o = n29605_o[2:0];
  /* ../../HW/src/dp/dp_gen.vhd:602:62  */
  assign n29805_o = n29803_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:603:42  */
  assign n29806_o = n29605_o[100:98];
  /* ../../HW/src/dp/dp_gen.vhd:603:62  */
  assign n29808_o = n29806_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:602:86  */
  assign n29809_o = n29808_o & n29805_o;
  /* ../../HW/src/dp/dp_gen.vhd:604:42  */
  assign n29810_o = n29605_o[198:196];
  /* ../../HW/src/dp/dp_gen.vhd:604:62  */
  assign n29812_o = n29810_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:603:86  */
  assign n29813_o = n29812_o & n29809_o;
  /* ../../HW/src/dp/dp_gen.vhd:605:42  */
  assign n29814_o = n29605_o[296:294];
  /* ../../HW/src/dp/dp_gen.vhd:605:62  */
  assign n29816_o = n29814_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:604:86  */
  assign n29817_o = n29816_o & n29813_o;
  /* ../../HW/src/dp/dp_gen.vhd:606:42  */
  assign n29818_o = n29605_o[394:392];
  /* ../../HW/src/dp/dp_gen.vhd:606:62  */
  assign n29820_o = n29818_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:605:86  */
  assign n29821_o = n29820_o & n29817_o;
  /* ../../HW/src/dp/dp_gen.vhd:607:35  */
  assign n29822_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:607:46  */
  assign n29824_o = n29822_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:606:86  */
  assign n29825_o = n29824_o & n29821_o;
  /* ../../HW/src/dp/dp_gen.vhd:608:40  */
  assign n29826_o = n29605_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:608:60  */
  assign n29828_o = n29826_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:607:105  */
  assign n29829_o = n29828_o & n29825_o;
  /* ../../HW/src/dp/dp_gen.vhd:609:44  */
  assign n29830_o = n29605_o[492:490];
  /* ../../HW/src/dp/dp_gen.vhd:609:64  */
  assign n29832_o = n29830_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:608:95  */
  assign n29833_o = n29832_o & n29829_o;
  /* ../../HW/src/dp/dp_gen.vhd:610:38  */
  assign n29834_o = n29605_o[595:593];
  /* ../../HW/src/dp/dp_gen.vhd:610:58  */
  assign n29836_o = n29834_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:609:99  */
  assign n29837_o = n29836_o & n29833_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:105  */
  assign n29838_o = n29802_o | n29837_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:5  */
  assign n29841_o = n29838_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:593:8  */
  assign n29842_o = n29785_o ? n29799_o : n29841_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:42  */
  assign n29843_o = n29604_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:541:62  */
  assign n29845_o = n29843_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:542:43  */
  assign n29847_o = pre_instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:541:98  */
  assign n29848_o = n29847_o & n29845_o;
  /* ../../HW/src/dp/dp_gen.vhd:543:37  */
  assign n29849_o = n29604_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:542:98  */
  assign n29850_o = n29849_o & n29848_o;
  /* ../../HW/src/dp/dp_gen.vhd:544:39  */
  assign n29851_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:544:50  */
  assign n29853_o = n29851_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:546:42  */
  assign n29854_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:546:53  */
  assign n29856_o = n29854_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:546:10  */
  assign n29857_o = n29856_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:544:10  */
  assign n29858_o = n29853_o ? 2'b01 : n29857_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:7  */
  assign n29859_o = n29850_o ? n29858_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:40  */
  assign n29860_o = n29605_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:555:60  */
  assign n29862_o = n29860_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:556:41  */
  assign n29864_o = pre_instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:96  */
  assign n29865_o = n29864_o & n29862_o;
  /* ../../HW/src/dp/dp_gen.vhd:557:35  */
  assign n29866_o = n29605_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:556:96  */
  assign n29867_o = n29866_o & n29865_o;
  /* ../../HW/src/dp/dp_gen.vhd:558:37  */
  assign n29868_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:558:48  */
  assign n29870_o = n29868_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:560:40  */
  assign n29871_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:560:51  */
  assign n29873_o = n29871_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:560:10  */
  assign n29874_o = n29873_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:558:10  */
  assign n29875_o = n29870_o ? 2'b01 : n29874_o;
  /* ../../HW/src/dp/dp_gen.vhd:555:7  */
  assign n29876_o = n29867_o ? n29875_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:569:42  */
  assign n29878_o = pre_instruction_bus_id_source_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:570:39  */
  assign n29879_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:570:50  */
  assign n29881_o = n29879_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:571:39  */
  assign n29882_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:571:50  */
  assign n29884_o = n29882_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:572:44  */
  assign n29885_o = n29604_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:572:64  */
  assign n29887_o = n29885_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:571:111  */
  assign n29888_o = n29887_o & n29884_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:111  */
  assign n29889_o = n29881_o | n29888_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:10  */
  assign n29892_o = n29889_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:577:39  */
  assign n29893_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:577:50  */
  assign n29895_o = n29893_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:578:46  */
  assign n29896_o = n29604_o[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:578:66  */
  assign n29898_o = n29896_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:579:46  */
  assign n29899_o = n29604_o[99:98];
  /* ../../HW/src/dp/dp_gen.vhd:579:66  */
  assign n29901_o = n29899_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:578:90  */
  assign n29902_o = n29901_o & n29898_o;
  /* ../../HW/src/dp/dp_gen.vhd:580:46  */
  assign n29903_o = n29604_o[197:196];
  /* ../../HW/src/dp/dp_gen.vhd:580:66  */
  assign n29905_o = n29903_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:579:90  */
  assign n29906_o = n29905_o & n29902_o;
  /* ../../HW/src/dp/dp_gen.vhd:581:46  */
  assign n29907_o = n29604_o[295:294];
  /* ../../HW/src/dp/dp_gen.vhd:581:66  */
  assign n29909_o = n29907_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:580:90  */
  assign n29910_o = n29909_o & n29906_o;
  /* ../../HW/src/dp/dp_gen.vhd:582:46  */
  assign n29911_o = n29604_o[393:392];
  /* ../../HW/src/dp/dp_gen.vhd:582:66  */
  assign n29913_o = n29911_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:581:90  */
  assign n29914_o = n29913_o & n29910_o;
  /* ../../HW/src/dp/dp_gen.vhd:583:39  */
  assign n29915_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:583:50  */
  assign n29917_o = n29915_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:582:90  */
  assign n29918_o = n29917_o & n29914_o;
  /* ../../HW/src/dp/dp_gen.vhd:584:44  */
  assign n29919_o = n29604_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:584:64  */
  assign n29921_o = n29919_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:583:111  */
  assign n29922_o = n29921_o & n29918_o;
  /* ../../HW/src/dp/dp_gen.vhd:585:48  */
  assign n29923_o = n29604_o[491:490];
  /* ../../HW/src/dp/dp_gen.vhd:585:68  */
  assign n29925_o = n29923_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:584:99  */
  assign n29926_o = n29925_o & n29922_o;
  /* ../../HW/src/dp/dp_gen.vhd:586:42  */
  assign n29927_o = n29604_o[594:593];
  /* ../../HW/src/dp/dp_gen.vhd:586:62  */
  assign n29929_o = n29927_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:585:103  */
  assign n29930_o = n29929_o & n29926_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:111  */
  assign n29931_o = n29895_o | n29930_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:7  */
  assign n29934_o = n29931_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:569:7  */
  assign n29935_o = n29878_o ? n29892_o : n29934_o;
  /* ../../HW/src/dp/dp_gen.vhd:593:41  */
  assign n29937_o = pre_instruction_bus_id_dest_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:594:38  */
  assign n29938_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:594:49  */
  assign n29940_o = n29938_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:595:38  */
  assign n29941_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:595:49  */
  assign n29943_o = n29941_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:596:43  */
  assign n29944_o = n29605_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:596:63  */
  assign n29946_o = n29944_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:595:108  */
  assign n29947_o = n29946_o & n29943_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:108  */
  assign n29948_o = n29940_o | n29947_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:11  */
  assign n29951_o = n29948_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:601:35  */
  assign n29952_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:601:46  */
  assign n29954_o = n29952_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:602:42  */
  assign n29955_o = n29605_o[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:602:62  */
  assign n29957_o = n29955_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:603:42  */
  assign n29958_o = n29605_o[99:98];
  /* ../../HW/src/dp/dp_gen.vhd:603:62  */
  assign n29960_o = n29958_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:602:86  */
  assign n29961_o = n29960_o & n29957_o;
  /* ../../HW/src/dp/dp_gen.vhd:604:42  */
  assign n29962_o = n29605_o[197:196];
  /* ../../HW/src/dp/dp_gen.vhd:604:62  */
  assign n29964_o = n29962_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:603:86  */
  assign n29965_o = n29964_o & n29961_o;
  /* ../../HW/src/dp/dp_gen.vhd:605:42  */
  assign n29966_o = n29605_o[295:294];
  /* ../../HW/src/dp/dp_gen.vhd:605:62  */
  assign n29968_o = n29966_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:604:86  */
  assign n29969_o = n29968_o & n29965_o;
  /* ../../HW/src/dp/dp_gen.vhd:606:42  */
  assign n29970_o = n29605_o[393:392];
  /* ../../HW/src/dp/dp_gen.vhd:606:62  */
  assign n29972_o = n29970_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:605:86  */
  assign n29973_o = n29972_o & n29969_o;
  /* ../../HW/src/dp/dp_gen.vhd:607:35  */
  assign n29974_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:607:46  */
  assign n29976_o = n29974_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:606:86  */
  assign n29977_o = n29976_o & n29973_o;
  /* ../../HW/src/dp/dp_gen.vhd:608:40  */
  assign n29978_o = n29605_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:608:60  */
  assign n29980_o = n29978_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:607:105  */
  assign n29981_o = n29980_o & n29977_o;
  /* ../../HW/src/dp/dp_gen.vhd:609:44  */
  assign n29982_o = n29605_o[491:490];
  /* ../../HW/src/dp/dp_gen.vhd:609:64  */
  assign n29984_o = n29982_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:608:95  */
  assign n29985_o = n29984_o & n29981_o;
  /* ../../HW/src/dp/dp_gen.vhd:610:38  */
  assign n29986_o = n29605_o[594:593];
  /* ../../HW/src/dp/dp_gen.vhd:610:58  */
  assign n29988_o = n29986_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:609:99  */
  assign n29989_o = n29988_o & n29985_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:105  */
  assign n29990_o = n29954_o | n29989_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:5  */
  assign n29993_o = n29990_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:593:8  */
  assign n29994_o = n29937_o ? n29951_o : n29993_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:42  */
  assign n29995_o = n29604_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:541:62  */
  assign n29997_o = n29995_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:542:43  */
  assign n29999_o = pre_instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:541:98  */
  assign n30000_o = n29999_o & n29997_o;
  /* ../../HW/src/dp/dp_gen.vhd:543:37  */
  assign n30001_o = n29604_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:542:98  */
  assign n30002_o = n30001_o & n30000_o;
  /* ../../HW/src/dp/dp_gen.vhd:544:39  */
  assign n30003_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:544:50  */
  assign n30005_o = n30003_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:546:42  */
  assign n30006_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:546:53  */
  assign n30008_o = n30006_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:546:10  */
  assign n30009_o = n30008_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:544:10  */
  assign n30010_o = n30005_o ? 2'b01 : n30009_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:7  */
  assign n30011_o = n30002_o ? n30010_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:40  */
  assign n30012_o = n29605_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:555:60  */
  assign n30014_o = n30012_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:556:41  */
  assign n30016_o = pre_instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:96  */
  assign n30017_o = n30016_o & n30014_o;
  /* ../../HW/src/dp/dp_gen.vhd:557:35  */
  assign n30018_o = n29605_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:556:96  */
  assign n30019_o = n30018_o & n30017_o;
  /* ../../HW/src/dp/dp_gen.vhd:558:37  */
  assign n30020_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:558:48  */
  assign n30022_o = n30020_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:560:40  */
  assign n30023_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:560:51  */
  assign n30025_o = n30023_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:560:10  */
  assign n30026_o = n30025_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:558:10  */
  assign n30027_o = n30022_o ? 2'b01 : n30026_o;
  /* ../../HW/src/dp/dp_gen.vhd:555:7  */
  assign n30028_o = n30019_o ? n30027_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:569:42  */
  assign n30030_o = pre_instruction_bus_id_source_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:570:39  */
  assign n30031_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:570:50  */
  assign n30033_o = n30031_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:571:39  */
  assign n30034_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:571:50  */
  assign n30036_o = n30034_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:572:44  */
  assign n30037_o = n29604_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:572:64  */
  assign n30039_o = n30037_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:571:111  */
  assign n30040_o = n30039_o & n30036_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:111  */
  assign n30041_o = n30033_o | n30040_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:10  */
  assign n30044_o = n30041_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:577:39  */
  assign n30045_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:577:50  */
  assign n30047_o = n30045_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:578:46  */
  assign n30048_o = n29604_o[0];
  /* ../../HW/src/dp/dp_gen.vhd:578:66  */
  assign n30050_o = n30048_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:579:46  */
  assign n30051_o = n29604_o[98];
  /* ../../HW/src/dp/dp_gen.vhd:579:66  */
  assign n30053_o = n30051_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:578:90  */
  assign n30054_o = n30053_o & n30050_o;
  /* ../../HW/src/dp/dp_gen.vhd:580:46  */
  assign n30055_o = n29604_o[196];
  /* ../../HW/src/dp/dp_gen.vhd:580:66  */
  assign n30057_o = n30055_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:579:90  */
  assign n30058_o = n30057_o & n30054_o;
  /* ../../HW/src/dp/dp_gen.vhd:581:46  */
  assign n30059_o = n29604_o[294];
  /* ../../HW/src/dp/dp_gen.vhd:581:66  */
  assign n30061_o = n30059_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:580:90  */
  assign n30062_o = n30061_o & n30058_o;
  /* ../../HW/src/dp/dp_gen.vhd:582:46  */
  assign n30063_o = n29604_o[392];
  /* ../../HW/src/dp/dp_gen.vhd:582:66  */
  assign n30065_o = n30063_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:581:90  */
  assign n30066_o = n30065_o & n30062_o;
  /* ../../HW/src/dp/dp_gen.vhd:583:39  */
  assign n30067_o = n29604_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:583:50  */
  assign n30069_o = n30067_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:582:90  */
  assign n30070_o = n30069_o & n30066_o;
  /* ../../HW/src/dp/dp_gen.vhd:584:44  */
  assign n30071_o = n29604_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:584:64  */
  assign n30073_o = n30071_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:583:111  */
  assign n30074_o = n30073_o & n30070_o;
  /* ../../HW/src/dp/dp_gen.vhd:585:48  */
  assign n30075_o = n29604_o[490];
  /* ../../HW/src/dp/dp_gen.vhd:585:68  */
  assign n30077_o = n30075_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:584:99  */
  assign n30078_o = n30077_o & n30074_o;
  /* ../../HW/src/dp/dp_gen.vhd:586:42  */
  assign n30079_o = n29604_o[593];
  /* ../../HW/src/dp/dp_gen.vhd:586:62  */
  assign n30081_o = n30079_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:585:103  */
  assign n30082_o = n30081_o & n30078_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:111  */
  assign n30083_o = n30047_o | n30082_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:7  */
  assign n30086_o = n30083_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:569:7  */
  assign n30087_o = n30030_o ? n30044_o : n30086_o;
  /* ../../HW/src/dp/dp_gen.vhd:593:41  */
  assign n30089_o = pre_instruction_bus_id_dest_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:594:38  */
  assign n30090_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:594:49  */
  assign n30092_o = n30090_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:595:38  */
  assign n30093_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:595:49  */
  assign n30095_o = n30093_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:596:43  */
  assign n30096_o = n29605_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:596:63  */
  assign n30098_o = n30096_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:595:108  */
  assign n30099_o = n30098_o & n30095_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:108  */
  assign n30100_o = n30092_o | n30099_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:11  */
  assign n30103_o = n30100_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:601:35  */
  assign n30104_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:601:46  */
  assign n30106_o = n30104_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:602:42  */
  assign n30107_o = n29605_o[0];
  /* ../../HW/src/dp/dp_gen.vhd:602:62  */
  assign n30109_o = n30107_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:603:42  */
  assign n30110_o = n29605_o[98];
  /* ../../HW/src/dp/dp_gen.vhd:603:62  */
  assign n30112_o = n30110_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:602:86  */
  assign n30113_o = n30112_o & n30109_o;
  /* ../../HW/src/dp/dp_gen.vhd:604:42  */
  assign n30114_o = n29605_o[196];
  /* ../../HW/src/dp/dp_gen.vhd:604:62  */
  assign n30116_o = n30114_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:603:86  */
  assign n30117_o = n30116_o & n30113_o;
  /* ../../HW/src/dp/dp_gen.vhd:605:42  */
  assign n30118_o = n29605_o[294];
  /* ../../HW/src/dp/dp_gen.vhd:605:62  */
  assign n30120_o = n30118_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:604:86  */
  assign n30121_o = n30120_o & n30117_o;
  /* ../../HW/src/dp/dp_gen.vhd:606:42  */
  assign n30122_o = n29605_o[392];
  /* ../../HW/src/dp/dp_gen.vhd:606:62  */
  assign n30124_o = n30122_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:605:86  */
  assign n30125_o = n30124_o & n30121_o;
  /* ../../HW/src/dp/dp_gen.vhd:607:35  */
  assign n30126_o = n29605_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:607:46  */
  assign n30128_o = n30126_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:606:86  */
  assign n30129_o = n30128_o & n30125_o;
  /* ../../HW/src/dp/dp_gen.vhd:608:40  */
  assign n30130_o = n29605_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:608:60  */
  assign n30132_o = n30130_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:607:105  */
  assign n30133_o = n30132_o & n30129_o;
  /* ../../HW/src/dp/dp_gen.vhd:609:44  */
  assign n30134_o = n29605_o[490];
  /* ../../HW/src/dp/dp_gen.vhd:609:64  */
  assign n30136_o = n30134_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:608:95  */
  assign n30137_o = n30136_o & n30133_o;
  /* ../../HW/src/dp/dp_gen.vhd:610:38  */
  assign n30138_o = n29605_o[593];
  /* ../../HW/src/dp/dp_gen.vhd:610:58  */
  assign n30140_o = n30138_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:609:99  */
  assign n30141_o = n30140_o & n30137_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:105  */
  assign n30142_o = n30106_o | n30141_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:5  */
  assign n30145_o = n30142_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:593:8  */
  assign n30146_o = n30089_o ? n30103_o : n30145_o;
  assign n30147_o = {n30087_o, n29935_o, n29783_o};
  assign n30149_o = {n30146_o, n29994_o, n29842_o};
  assign n30151_o = {n30011_o, n29859_o, n29707_o};
  assign n30153_o = {n30028_o, n29876_o, n29724_o};
  /* ../../HW/src/dp/dp_gen.vhd:627:21  */
  assign n30172_o = src_is_vector_r[0];
  /* ../../HW/src/dp/dp_gen.vhd:627:48  */
  assign n30173_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:627:51  */
  assign n30175_o = n30173_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:627:29  */
  assign n30176_o = n30172_o | n30175_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:95  */
  assign n30177_o = n29602_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:627:111  */
  assign n30178_o = ~n30177_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:69  */
  assign n30179_o = n30178_o & n30176_o;
  /* ../../HW/src/dp/dp_gen.vhd:628:21  */
  assign n30180_o = dst_is_vector_r[0];
  /* ../../HW/src/dp/dp_gen.vhd:628:48  */
  assign n30181_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:628:51  */
  assign n30183_o = n30181_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:628:29  */
  assign n30184_o = n30180_o | n30183_o;
  /* ../../HW/src/dp/dp_gen.vhd:628:93  */
  assign n30185_o = n29603_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:628:109  */
  assign n30186_o = ~n30185_o;
  /* ../../HW/src/dp/dp_gen.vhd:628:69  */
  assign n30187_o = n30186_o & n30184_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:117  */
  assign n30188_o = n30187_o & n30179_o;
  /* ../../HW/src/dp/dp_gen.vhd:631:35  */
  assign n30189_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:632:35  */
  assign n30190_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:633:23  */
  assign n30191_o = src_is_vector_r[1];
  /* ../../HW/src/dp/dp_gen.vhd:633:50  */
  assign n30192_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:633:53  */
  assign n30194_o = n30192_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:633:31  */
  assign n30195_o = n30191_o | n30194_o;
  /* ../../HW/src/dp/dp_gen.vhd:634:23  */
  assign n30196_o = dst_is_vector_r[1];
  /* ../../HW/src/dp/dp_gen.vhd:634:50  */
  assign n30197_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:634:53  */
  assign n30199_o = n30197_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:634:31  */
  assign n30200_o = n30196_o | n30199_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:71  */
  assign n30201_o = n30200_o & n30195_o;
  /* ../../HW/src/dp/dp_gen.vhd:637:35  */
  assign n30202_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:638:35  */
  assign n30203_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:639:23  */
  assign n30204_o = src_is_vector_r[2];
  /* ../../HW/src/dp/dp_gen.vhd:639:50  */
  assign n30205_o = src_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:639:53  */
  assign n30207_o = n30205_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:639:31  */
  assign n30208_o = n30204_o | n30207_o;
  /* ../../HW/src/dp/dp_gen.vhd:640:23  */
  assign n30209_o = dst_is_vector_r[2];
  /* ../../HW/src/dp/dp_gen.vhd:640:50  */
  assign n30210_o = dst_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:640:53  */
  assign n30212_o = n30210_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:640:31  */
  assign n30213_o = n30209_o | n30212_o;
  /* ../../HW/src/dp/dp_gen.vhd:639:71  */
  assign n30214_o = n30213_o & n30208_o;
  /* ../../HW/src/dp/dp_gen.vhd:643:35  */
  assign n30215_o = src_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:644:35  */
  assign n30216_o = dst_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n30219_o = n30214_o ? 3'b001 : 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n30222_o = n30214_o ? 3'b001 : 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n30224_o = n30214_o ? n30215_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n30226_o = n30214_o ? n30216_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n30228_o = n30201_o ? 3'b011 : n30219_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n30230_o = n30201_o ? 3'b011 : n30222_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n30231_o = n30201_o ? n30202_o : n30224_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n30232_o = n30201_o ? n30203_o : n30226_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n30234_o = n30188_o ? 3'b111 : n30228_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n30236_o = n30188_o ? 3'b111 : n30230_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n30237_o = n30188_o ? n30189_o : n30231_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n30238_o = n30188_o ? n30190_o : n30232_o;
  /* ../../HW/src/dp/dp_gen.vhd:658:31  */
  assign n30241_o = s_burstlen_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:659:56  */
  assign n30242_o = s_template_r[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:659:31  */
  assign n30243_o = s_burstpos_r + n30242_o;
  /* ../../HW/src/dp/dp_gen.vhd:660:40  */
  assign n30244_o = s_template_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:660:19  */
  assign n30245_o = s_i0_r + n30244_o;
  /* ../../HW/src/dp/dp_gen.vhd:661:40  */
  assign n30246_o = s_template_r[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:661:19  */
  assign n30247_o = s_i1_r + n30246_o;
  /* ../../HW/src/dp/dp_gen.vhd:662:40  */
  assign n30248_o = s_template_r[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:662:19  */
  assign n30249_o = s_i2_r + n30248_o;
  /* ../../HW/src/dp/dp_gen.vhd:663:40  */
  assign n30250_o = s_template_r[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:663:19  */
  assign n30251_o = s_i3_r + n30250_o;
  /* ../../HW/src/dp/dp_gen.vhd:664:40  */
  assign n30252_o = s_template_r[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:664:19  */
  assign n30253_o = s_i4_r + n30252_o;
  /* ../../HW/src/dp/dp_gen.vhd:666:57  */
  assign n30255_o = {1'b0, s_burstpos_stride_r};
  /* ../../HW/src/dp/dp_gen.vhd:666:43  */
  assign n30256_o = s_burstpos_start_r + n30255_o;
  /* ../../HW/src/dp/dp_gen.vhd:667:84  */
  assign n30257_o = s_template_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:667:45  */
  assign n30259_o = {1'b0, n30257_o};
  /* ../../HW/src/dp/dp_gen.vhd:667:31  */
  assign n30260_o = s_i0_start_r + n30259_o;
  /* ../../HW/src/dp/dp_gen.vhd:668:84  */
  assign n30261_o = s_template_r[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:668:45  */
  assign n30263_o = {1'b0, n30261_o};
  /* ../../HW/src/dp/dp_gen.vhd:668:31  */
  assign n30264_o = s_i1_start_r + n30263_o;
  /* ../../HW/src/dp/dp_gen.vhd:669:84  */
  assign n30265_o = s_template_r[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:669:45  */
  assign n30267_o = {1'b0, n30265_o};
  /* ../../HW/src/dp/dp_gen.vhd:669:31  */
  assign n30268_o = s_i2_start_r + n30267_o;
  /* ../../HW/src/dp/dp_gen.vhd:670:84  */
  assign n30269_o = s_template_r[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:670:45  */
  assign n30271_o = {1'b0, n30269_o};
  /* ../../HW/src/dp/dp_gen.vhd:670:31  */
  assign n30272_o = s_i3_start_r + n30271_o;
  /* ../../HW/src/dp/dp_gen.vhd:671:84  */
  assign n30273_o = s_template_r[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:671:45  */
  assign n30275_o = {1'b0, n30273_o};
  /* ../../HW/src/dp/dp_gen.vhd:671:31  */
  assign n30276_o = s_i4_start_r + n30275_o;
  /* ../../HW/src/dp/dp_gen.vhd:673:31  */
  assign n30278_o = s_i0_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:674:31  */
  assign n30280_o = s_i1_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:675:31  */
  assign n30282_o = s_i2_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:676:31  */
  assign n30284_o = s_i3_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:677:31  */
  assign n30286_o = s_i4_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:679:31  */
  assign n30288_o = d_burstlen_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:680:45  */
  assign n30289_o = d_template_r[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:680:31  */
  assign n30290_o = d_burstpos_r + n30289_o;
  /* ../../HW/src/dp/dp_gen.vhd:681:33  */
  assign n30291_o = d_template_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:681:19  */
  assign n30292_o = d_i0_r + n30291_o;
  /* ../../HW/src/dp/dp_gen.vhd:682:33  */
  assign n30293_o = d_template_r[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:682:19  */
  assign n30294_o = d_i1_r + n30293_o;
  /* ../../HW/src/dp/dp_gen.vhd:683:33  */
  assign n30295_o = d_template_r[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:683:19  */
  assign n30296_o = d_i2_r + n30295_o;
  /* ../../HW/src/dp/dp_gen.vhd:684:33  */
  assign n30297_o = d_template_r[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:684:19  */
  assign n30298_o = d_i3_r + n30297_o;
  /* ../../HW/src/dp/dp_gen.vhd:685:33  */
  assign n30299_o = d_template_r[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:685:19  */
  assign n30300_o = d_i4_r + n30299_o;
  /* ../../HW/src/dp/dp_gen.vhd:687:68  */
  assign n30301_o = d_template_r[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:687:97  */
  assign n30303_o = {n30301_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:687:20  */
  assign n30304_o = d_i0_r + n30303_o;
  /* ../../HW/src/dp/dp_gen.vhd:688:68  */
  assign n30305_o = d_template_r[120:98];
  /* ../../HW/src/dp/dp_gen.vhd:688:97  */
  assign n30307_o = {n30305_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:688:20  */
  assign n30308_o = d_i1_r + n30307_o;
  /* ../../HW/src/dp/dp_gen.vhd:689:68  */
  assign n30309_o = d_template_r[218:196];
  /* ../../HW/src/dp/dp_gen.vhd:689:97  */
  assign n30311_o = {n30309_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:689:20  */
  assign n30312_o = d_i2_r + n30311_o;
  /* ../../HW/src/dp/dp_gen.vhd:690:68  */
  assign n30313_o = d_template_r[316:294];
  /* ../../HW/src/dp/dp_gen.vhd:690:97  */
  assign n30315_o = {n30313_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:690:20  */
  assign n30316_o = d_i3_r + n30315_o;
  /* ../../HW/src/dp/dp_gen.vhd:691:68  */
  assign n30317_o = d_template_r[414:392];
  /* ../../HW/src/dp/dp_gen.vhd:691:97  */
  assign n30319_o = {n30317_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:691:20  */
  assign n30320_o = d_i4_r + n30319_o;
  /* ../../HW/src/dp/dp_gen.vhd:693:31  */
  assign n30322_o = d_i0_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:694:31  */
  assign n30324_o = d_i1_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:695:31  */
  assign n30326_o = d_i2_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:696:31  */
  assign n30328_o = d_i3_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:697:31  */
  assign n30330_o = d_i4_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:712:67  */
  assign n30333_o = ~s_gen_burstlen_progress_r;
  /* ../../HW/src/dp/dp_gen.vhd:712:39  */
  assign n30334_o = eof_rrrr | n30333_o;
  /* ../../HW/src/dp/dp_gen.vhd:712:20  */
  assign n30335_o = n30334_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:719:33  */
  assign n30338_o = waitreq_in & gen_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:719:49  */
  assign n30340_o = n30338_o != 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:719:16  */
  assign n30341_o = n30340_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:725:82  */
  assign n30344_o = s_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:725:53  */
  assign n30345_o = s_burstlen_r == n30344_o;
  /* ../../HW/src/dp/dp_gen.vhd:725:24  */
  assign n30346_o = n30345_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:726:84  */
  assign n30349_o = s_template_r[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:726:47  */
  assign n30350_o = s_i0_count_r == n30349_o;
  /* ../../HW/src/dp/dp_gen.vhd:726:18  */
  assign n30351_o = n30350_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:727:84  */
  assign n30354_o = s_template_r[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:727:47  */
  assign n30355_o = s_i1_count_r == n30354_o;
  /* ../../HW/src/dp/dp_gen.vhd:727:18  */
  assign n30356_o = n30355_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:728:84  */
  assign n30359_o = s_template_r[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:728:47  */
  assign n30360_o = s_i2_count_r == n30359_o;
  /* ../../HW/src/dp/dp_gen.vhd:728:18  */
  assign n30361_o = n30360_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:729:84  */
  assign n30364_o = s_template_r[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:729:47  */
  assign n30365_o = s_i3_count_r == n30364_o;
  /* ../../HW/src/dp/dp_gen.vhd:729:18  */
  assign n30366_o = n30365_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:730:84  */
  assign n30369_o = s_template_r[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:730:47  */
  assign n30370_o = s_i4_count_r == n30369_o;
  /* ../../HW/src/dp/dp_gen.vhd:730:18  */
  assign n30371_o = n30370_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:732:78  */
  assign n30374_o = s_template_r[71:48];
  /* ../../HW/src/dp/dp_gen.vhd:732:42  */
  assign n30375_o = $unsigned(s_i0_r) <= $unsigned(n30374_o);
  /* ../../HW/src/dp/dp_gen.vhd:732:136  */
  assign n30376_o = s_template_r[72];
  /* ../../HW/src/dp/dp_gen.vhd:732:153  */
  assign n30377_o = ~n30376_o;
  /* ../../HW/src/dp/dp_gen.vhd:732:108  */
  assign n30378_o = n30377_o & n30375_o;
  /* ../../HW/src/dp/dp_gen.vhd:732:19  */
  assign n30379_o = n30378_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:733:78  */
  assign n30382_o = s_template_r[169:146];
  /* ../../HW/src/dp/dp_gen.vhd:733:42  */
  assign n30383_o = $unsigned(s_i1_r) <= $unsigned(n30382_o);
  /* ../../HW/src/dp/dp_gen.vhd:733:136  */
  assign n30384_o = s_template_r[170];
  /* ../../HW/src/dp/dp_gen.vhd:733:153  */
  assign n30385_o = ~n30384_o;
  /* ../../HW/src/dp/dp_gen.vhd:733:108  */
  assign n30386_o = n30385_o & n30383_o;
  /* ../../HW/src/dp/dp_gen.vhd:733:19  */
  assign n30387_o = n30386_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:734:78  */
  assign n30390_o = s_template_r[267:244];
  /* ../../HW/src/dp/dp_gen.vhd:734:42  */
  assign n30391_o = $unsigned(s_i2_r) <= $unsigned(n30390_o);
  /* ../../HW/src/dp/dp_gen.vhd:734:136  */
  assign n30392_o = s_template_r[268];
  /* ../../HW/src/dp/dp_gen.vhd:734:153  */
  assign n30393_o = ~n30392_o;
  /* ../../HW/src/dp/dp_gen.vhd:734:108  */
  assign n30394_o = n30393_o & n30391_o;
  /* ../../HW/src/dp/dp_gen.vhd:734:19  */
  assign n30395_o = n30394_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:735:78  */
  assign n30398_o = s_template_r[365:342];
  /* ../../HW/src/dp/dp_gen.vhd:735:42  */
  assign n30399_o = $unsigned(s_i3_r) <= $unsigned(n30398_o);
  /* ../../HW/src/dp/dp_gen.vhd:735:136  */
  assign n30400_o = s_template_r[366];
  /* ../../HW/src/dp/dp_gen.vhd:735:153  */
  assign n30401_o = ~n30400_o;
  /* ../../HW/src/dp/dp_gen.vhd:735:108  */
  assign n30402_o = n30401_o & n30399_o;
  /* ../../HW/src/dp/dp_gen.vhd:735:19  */
  assign n30403_o = n30402_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:736:78  */
  assign n30406_o = s_template_r[463:440];
  /* ../../HW/src/dp/dp_gen.vhd:736:42  */
  assign n30407_o = $unsigned(s_i4_r) <= $unsigned(n30406_o);
  /* ../../HW/src/dp/dp_gen.vhd:736:136  */
  assign n30408_o = s_template_r[464];
  /* ../../HW/src/dp/dp_gen.vhd:736:153  */
  assign n30409_o = ~n30408_o;
  /* ../../HW/src/dp/dp_gen.vhd:736:108  */
  assign n30410_o = n30409_o & n30407_o;
  /* ../../HW/src/dp/dp_gen.vhd:736:19  */
  assign n30411_o = n30410_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:737:85  */
  assign n30414_o = s_template_r[513:490];
  /* ../../HW/src/dp/dp_gen.vhd:737:51  */
  assign n30415_o = $unsigned(s_burstpos_r) <= $unsigned(n30414_o);
  /* ../../HW/src/dp/dp_gen.vhd:737:141  */
  assign n30416_o = s_template_r[514];
  /* ../../HW/src/dp/dp_gen.vhd:737:158  */
  assign n30417_o = ~n30416_o;
  /* ../../HW/src/dp/dp_gen.vhd:737:115  */
  assign n30418_o = n30417_o & n30415_o;
  /* ../../HW/src/dp/dp_gen.vhd:737:22  */
  assign n30419_o = n30418_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:739:37  */
  assign n30421_o = s_i0_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:739:21  */
  assign n30422_o = ~n30421_o;
  /* ../../HW/src/dp/dp_gen.vhd:740:37  */
  assign n30423_o = s_i1_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:740:21  */
  assign n30424_o = ~n30423_o;
  /* ../../HW/src/dp/dp_gen.vhd:741:37  */
  assign n30425_o = s_i2_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:741:21  */
  assign n30426_o = ~n30425_o;
  /* ../../HW/src/dp/dp_gen.vhd:742:37  */
  assign n30427_o = s_i3_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:742:21  */
  assign n30428_o = ~n30427_o;
  /* ../../HW/src/dp/dp_gen.vhd:743:37  */
  assign n30429_o = s_i4_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:743:21  */
  assign n30430_o = ~n30429_o;
  /* ../../HW/src/dp/dp_gen.vhd:744:61  */
  assign n30432_o = {{1{s_burstpos_stride_r[23]}}, s_burstpos_stride_r}; // sext
  /* ../../HW/src/dp/dp_gen.vhd:744:61  */
  assign n30433_o = s_burstpos_start_r + n30432_o;
  /* ../../HW/src/dp/dp_gen.vhd:744:91  */
  assign n30435_o = $signed(n30433_o) >= $signed(25'b0000000000000000000000001);
  /* ../../HW/src/dp/dp_gen.vhd:744:28  */
  assign n30436_o = n30435_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:746:77  */
  assign n30439_o = d_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:746:53  */
  assign n30440_o = d_burstlen_r == n30439_o;
  /* ../../HW/src/dp/dp_gen.vhd:746:24  */
  assign n30441_o = n30440_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:747:71  */
  assign n30444_o = d_template_r[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:747:47  */
  assign n30445_o = d_i0_count_r == n30444_o;
  /* ../../HW/src/dp/dp_gen.vhd:747:18  */
  assign n30446_o = n30445_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:748:71  */
  assign n30449_o = d_template_r[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:748:47  */
  assign n30450_o = d_i1_count_r == n30449_o;
  /* ../../HW/src/dp/dp_gen.vhd:748:18  */
  assign n30451_o = n30450_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:749:71  */
  assign n30454_o = d_template_r[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:749:47  */
  assign n30455_o = d_i2_count_r == n30454_o;
  /* ../../HW/src/dp/dp_gen.vhd:749:18  */
  assign n30456_o = n30455_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:750:71  */
  assign n30459_o = d_template_r[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:750:47  */
  assign n30460_o = d_i3_count_r == n30459_o;
  /* ../../HW/src/dp/dp_gen.vhd:750:18  */
  assign n30461_o = n30460_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:751:71  */
  assign n30464_o = d_template_r[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:751:47  */
  assign n30465_o = d_i4_count_r == n30464_o;
  /* ../../HW/src/dp/dp_gen.vhd:751:18  */
  assign n30466_o = n30465_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:753:78  */
  assign n30469_o = d_template_r[71:48];
  /* ../../HW/src/dp/dp_gen.vhd:753:42  */
  assign n30470_o = $unsigned(d_i0_r) <= $unsigned(n30469_o);
  /* ../../HW/src/dp/dp_gen.vhd:753:136  */
  assign n30471_o = d_template_r[72];
  /* ../../HW/src/dp/dp_gen.vhd:753:153  */
  assign n30472_o = ~n30471_o;
  /* ../../HW/src/dp/dp_gen.vhd:753:108  */
  assign n30473_o = n30472_o & n30470_o;
  /* ../../HW/src/dp/dp_gen.vhd:753:19  */
  assign n30474_o = n30473_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:754:78  */
  assign n30477_o = d_template_r[169:146];
  /* ../../HW/src/dp/dp_gen.vhd:754:42  */
  assign n30478_o = $unsigned(d_i1_r) <= $unsigned(n30477_o);
  /* ../../HW/src/dp/dp_gen.vhd:754:136  */
  assign n30479_o = d_template_r[170];
  /* ../../HW/src/dp/dp_gen.vhd:754:153  */
  assign n30480_o = ~n30479_o;
  /* ../../HW/src/dp/dp_gen.vhd:754:108  */
  assign n30481_o = n30480_o & n30478_o;
  /* ../../HW/src/dp/dp_gen.vhd:754:19  */
  assign n30482_o = n30481_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:755:78  */
  assign n30485_o = d_template_r[267:244];
  /* ../../HW/src/dp/dp_gen.vhd:755:42  */
  assign n30486_o = $unsigned(d_i2_r) <= $unsigned(n30485_o);
  /* ../../HW/src/dp/dp_gen.vhd:755:136  */
  assign n30487_o = d_template_r[268];
  /* ../../HW/src/dp/dp_gen.vhd:755:153  */
  assign n30488_o = ~n30487_o;
  /* ../../HW/src/dp/dp_gen.vhd:755:108  */
  assign n30489_o = n30488_o & n30486_o;
  /* ../../HW/src/dp/dp_gen.vhd:755:19  */
  assign n30490_o = n30489_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:756:78  */
  assign n30493_o = d_template_r[365:342];
  /* ../../HW/src/dp/dp_gen.vhd:756:42  */
  assign n30494_o = $unsigned(d_i3_r) <= $unsigned(n30493_o);
  /* ../../HW/src/dp/dp_gen.vhd:756:136  */
  assign n30495_o = d_template_r[366];
  /* ../../HW/src/dp/dp_gen.vhd:756:153  */
  assign n30496_o = ~n30495_o;
  /* ../../HW/src/dp/dp_gen.vhd:756:108  */
  assign n30497_o = n30496_o & n30494_o;
  /* ../../HW/src/dp/dp_gen.vhd:756:19  */
  assign n30498_o = n30497_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:757:78  */
  assign n30501_o = d_template_r[463:440];
  /* ../../HW/src/dp/dp_gen.vhd:757:42  */
  assign n30502_o = $unsigned(d_i4_r) <= $unsigned(n30501_o);
  /* ../../HW/src/dp/dp_gen.vhd:757:136  */
  assign n30503_o = d_template_r[464];
  /* ../../HW/src/dp/dp_gen.vhd:757:153  */
  assign n30504_o = ~n30503_o;
  /* ../../HW/src/dp/dp_gen.vhd:757:108  */
  assign n30505_o = n30504_o & n30502_o;
  /* ../../HW/src/dp/dp_gen.vhd:757:19  */
  assign n30506_o = n30505_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:758:76  */
  assign n30509_o = d_burst_max_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:758:51  */
  assign n30510_o = $unsigned(d_burstpos_r) <= $unsigned(n30509_o);
  /* ../../HW/src/dp/dp_gen.vhd:758:123  */
  assign n30511_o = d_burst_max_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:758:140  */
  assign n30512_o = ~n30511_o;
  /* ../../HW/src/dp/dp_gen.vhd:758:106  */
  assign n30513_o = n30512_o & n30510_o;
  /* ../../HW/src/dp/dp_gen.vhd:758:22  */
  assign n30514_o = n30513_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:776:16  */
  assign n30526_o = ~reset_in;
  /* ../../HW/src/dp/dp_gen.vhd:915:24  */
  assign n30528_o = ~waitreq;
  /* ../../HW/src/dp/dp_gen.vhd:920:40  */
  assign n30530_o = dp_src_bus_id_rrr == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:920:20  */
  assign n30532_o = n30530_o ? running_rrr : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:920:40  */
  assign n30534_o = dp_src_bus_id_rrr == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:920:20  */
  assign n30536_o = n30534_o ? running_rrr : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:920:40  */
  assign n30538_o = dp_src_bus_id_rrr == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:920:20  */
  assign n30540_o = n30538_o ? running_rrr : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:971:36  */
  assign n30544_o = s_i0_r + s_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:971:43  */
  assign n30545_o = n30544_o + s_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:972:52  */
  assign n30546_o = s_template_r[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:974:46  */
  assign n30547_o = s_template_r[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:975:48  */
  assign n30548_o = s_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:975:76  */
  assign n30549_o = n30548_o - s_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:976:42  */
  assign n30550_o = s_burstpos_r + s_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:976:49  */
  assign n30551_o = n30550_o + s_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:977:39  */
  assign n30552_o = s_temp1_r + s_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:979:27  */
  assign n30553_o = {8'b0, s_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:979:75  */
  assign n30554_o = n30553_o + s_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:981:43  */
  assign n30556_o = n30554_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:980:17  */
  assign n30557_o = src_double_rrr ? n30556_o : n30554_o;
  /* ../../HW/src/dp/dp_gen.vhd:985:37  */
  assign n30561_o = $unsigned(s_gen_burstlen_r) > $unsigned(n32878_o);
  /* ../../HW/src/dp/dp_gen.vhd:985:17  */
  assign n30565_o = n30561_o ? n32885_o : s_gen_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:991:34  */
  assign n30567_o = n30565_o == 5'b00000;
  /* ../../HW/src/dp/dp_gen.vhd:991:17  */
  assign n30570_o = n30567_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:1001:40  */
  assign n30571_o = {3'b0, s_burstpos_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1002:65  */
  assign n30572_o = s_burst_actual_max_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1002:38  */
  assign n30573_o = {3'b0, n30572_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1002:110  */
  assign n30574_o = n30573_o - n30571_o;
  /* ../../HW/src/dp/dp_gen.vhd:1002:122  */
  assign n30576_o = n30574_o + 27'b000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1004:39  */
  assign n30578_o = n30576_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1003:17  */
  assign n30579_o = src_double_r ? n30578_o : n30576_o;
  /* ../../HW/src/dp/dp_gen.vhd:1007:36  */
  assign n30580_o = s_burstpos_end_r[26];
  /* ../../HW/src/dp/dp_gen.vhd:1010:39  */
  assign n30581_o = s_burstpos_end_r[26:4];
  /* ../../HW/src/dp/dp_gen.vhd:1010:94  */
  assign n30583_o = n30581_o == 23'b00000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1012:57  */
  assign n30584_o = s_burstpos_end_r[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1010:17  */
  assign n30586_o = n30583_o ? n30584_o : 4'b1111;
  /* ../../HW/src/dp/dp_gen.vhd:1007:17  */
  assign n30588_o = n30580_o ? 4'b0000 : n30586_o;
  /* ../../HW/src/dp/dp_gen.vhd:1020:55  */
  assign n30589_o = s_bufsize_rr[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:1020:36  */
  assign n30590_o = {2'b0, n30589_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1020:111  */
  assign n30591_o = {1'b0, s_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1020:103  */
  assign n30592_o = n30590_o - n30591_o;
  /* ../../HW/src/dp/dp_gen.vhd:1022:41  */
  assign n30594_o = n30592_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1021:17  */
  assign n30595_o = src_double_rrr ? n30594_o : n30592_o;
  /* ../../HW/src/dp/dp_gen.vhd:1024:29  */
  assign n30597_o = $signed(n30595_o) <= $signed(25'b0000000000000000000000000);
  /* ../../HW/src/dp/dp_gen.vhd:1026:44  */
  assign n30598_o = {21'b0, s_burstpos_end_rr};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1026:42  */
  assign n30599_o = $unsigned(n30595_o) > $unsigned(n30598_o);
  /* ../../HW/src/dp/dp_gen.vhd:1029:59  */
  assign n30600_o = n30595_o[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1026:17  */
  assign n30601_o = n30599_o ? s_burstpos_end_rr : n30600_o;
  /* ../../HW/src/dp/dp_gen.vhd:1024:17  */
  assign n30603_o = n30597_o ? 4'b0000 : n30601_o;
  /* ../../HW/src/dp/dp_gen.vhd:1032:89  */
  assign n30605_o = s_template_r[512:490];
  /* ../../HW/src/dp/dp_gen.vhd:1032:47  */
  assign n30607_o = {1'b0, n30605_o};
  /* ../../HW/src/dp/dp_gen.vhd:1032:120  */
  assign n30608_o = n30607_o - s_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1033:42  */
  assign n30610_o = src_vector_r == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1034:106  */
  assign n30611_o = n30608_o[23:1];
  /* ../../HW/src/dp/dp_gen.vhd:1036:45  */
  assign n30614_o = src_vector_r == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1037:106  */
  assign n30615_o = n30608_o[23:2];
  /* ../../HW/src/dp/dp_gen.vhd:1039:45  */
  assign n30618_o = src_vector_r == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1040:104  */
  assign n30619_o = n30608_o[23:3];
  assign n30621_o = {3'b000, n30619_o};
  /* ../../HW/src/dp/dp_gen.vhd:1039:17  */
  assign n30622_o = n30618_o ? n30621_o : n30608_o;
  assign n30623_o = {2'b00, n30615_o};
  /* ../../HW/src/dp/dp_gen.vhd:1036:17  */
  assign n30624_o = n30614_o ? n30623_o : n30622_o;
  assign n30625_o = {1'b0, n30611_o};
  /* ../../HW/src/dp/dp_gen.vhd:1033:17  */
  assign n30626_o = n30610_o ? n30625_o : n30624_o;
  /* ../../HW/src/dp/dp_gen.vhd:1045:42  */
  assign n30627_o = s_i0_valid & s_i1_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:57  */
  assign n30628_o = n30627_o & s_i2_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:72  */
  assign n30629_o = n30628_o & s_i3_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:87  */
  assign n30630_o = n30629_o & s_i4_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:102  */
  assign n30631_o = n30630_o & s_burst_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:48  */
  assign n30632_o = s_i0_start_valid & s_i1_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:69  */
  assign n30633_o = n30632_o & s_i2_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:90  */
  assign n30634_o = n30633_o & s_i3_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:111  */
  assign n30635_o = n30634_o & s_i4_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:132  */
  assign n30636_o = n30635_o & s_burst_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:121  */
  assign n30637_o = n30631_o & n30636_o;
  /* ../../HW/src/dp/dp_gen.vhd:1047:29  */
  assign n30638_o = ~s_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:1049:45  */
  assign n30640_o = src_is_burst_rr & 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:1050:33  */
  assign n30641_o = s_temp3_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1050:78  */
  assign n30643_o = n30641_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1051:32  */
  assign n30644_o = s_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1051:62  */
  assign n30646_o = n30644_o != 5'b11111;
  /* ../../HW/src/dp/dp_gen.vhd:1050:129  */
  assign n30647_o = n30646_o & n30643_o;
  /* ../../HW/src/dp/dp_gen.vhd:1052:48  */
  assign n30648_o = s_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1050:20  */
  assign n30650_o = n30647_o ? n30648_o : 5'b11110;
  /* ../../HW/src/dp/dp_gen.vhd:1056:38  */
  assign n30651_o = s_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1058:41  */
  assign n30652_o = s_burstremain_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1058:92  */
  assign n30654_o = n30652_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1059:53  */
  assign n30655_o = s_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1059:36  */
  assign n30656_o = $unsigned(n30650_o) > $unsigned(n30655_o);
  /* ../../HW/src/dp/dp_gen.vhd:1058:149  */
  assign n30657_o = n30656_o & n30654_o;
  /* ../../HW/src/dp/dp_gen.vhd:1060:58  */
  assign n30658_o = s_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1060:88  */
  assign n30660_o = n30658_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1062:55  */
  assign n30662_o = n30650_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1058:20  */
  assign n30663_o = n30657_o ? n30660_o : n30662_o;
  /* ../../HW/src/dp/dp_gen.vhd:1056:20  */
  assign n30665_o = n30651_o ? 5'b00000 : n30663_o;
  /* ../../HW/src/dp/dp_gen.vhd:1065:38  */
  assign n30666_o = s_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1065:20  */
  assign n30669_o = n30666_o ? 5'b00000 : 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1049:17  */
  assign n30670_o = n30640_o ? n30665_o : n30669_o;
  /* ../../HW/src/dp/dp_gen.vhd:1047:17  */
  assign n30673_o = n30638_o ? 5'b00000 : n30670_o;
  /* ../../HW/src/dp/dp_gen.vhd:1103:84  */
  assign n30675_o = src_vector_rrr[1:0];
  assign n30677_o = {n30675_o, 1'b1};
  /* ../../HW/src/dp/dp_gen.vhd:1102:17  */
  assign n30678_o = src_double_rrr ? n30677_o : src_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:1112:38  */
  assign n30679_o = s_burstpos_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:1112:67  */
  assign n30680_o = ~n30679_o;
  /* ../../HW/src/dp/dp_gen.vhd:1115:41  */
  assign n30681_o = s_burstpos_start_r[24:3];
  /* ../../HW/src/dp/dp_gen.vhd:1115:96  */
  assign n30683_o = n30681_o == 22'b1111111111111111111111;
  /* ../../HW/src/dp/dp_gen.vhd:1117:61  */
  assign n30684_o = s_burstpos_start_r[3:0];
  assign n30687_o = {1'b1, 3'b000};
  /* ../../HW/src/dp/dp_gen.vhd:1115:17  */
  assign n30688_o = n30683_o ? n30684_o : n30687_o;
  /* ../../HW/src/dp/dp_gen.vhd:1112:17  */
  assign n30690_o = n30680_o ? 4'b0000 : n30688_o;
  /* ../../HW/src/dp/dp_gen.vhd:1129:84  */
  assign n30691_o = dst_vector_rrr[1:0];
  assign n30693_o = {n30691_o, 1'b1};
  /* ../../HW/src/dp/dp_gen.vhd:1128:17  */
  assign n30694_o = dst_double_rrr ? n30693_o : dst_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:1155:52  */
  assign n30695_o = d_template_r[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:1157:36  */
  assign n30696_o = d_i0_r + d_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:1157:43  */
  assign n30697_o = n30696_o + d_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:1158:43  */
  assign n30698_o = d_template_r[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:1159:43  */
  assign n30699_o = d_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:1159:48  */
  assign n30700_o = n30699_o - d_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1160:42  */
  assign n30701_o = d_burstpos_r + d_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:1160:49  */
  assign n30702_o = n30701_o + d_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1161:39  */
  assign n30703_o = d_temp1_r + d_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1164:27  */
  assign n30704_o = {8'b0, d_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1164:75  */
  assign n30705_o = n30704_o + d_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:1166:43  */
  assign n30707_o = n30705_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1165:17  */
  assign n30708_o = dst_double_rrr ? n30707_o : n30705_o;
  /* ../../HW/src/dp/dp_gen.vhd:1173:40  */
  assign n30709_o = {3'b0, d_burstpos_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1174:58  */
  assign n30710_o = d_burst_max_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1174:38  */
  assign n30711_o = {3'b0, n30710_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1174:103  */
  assign n30712_o = n30711_o - n30709_o;
  /* ../../HW/src/dp/dp_gen.vhd:1174:115  */
  assign n30714_o = n30712_o + 27'b000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1176:39  */
  assign n30716_o = n30714_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1175:17  */
  assign n30717_o = dst_double_r ? n30716_o : n30714_o;
  /* ../../HW/src/dp/dp_gen.vhd:1179:36  */
  assign n30718_o = d_burstpos_end_r[26];
  /* ../../HW/src/dp/dp_gen.vhd:1181:39  */
  assign n30719_o = d_burstpos_end_r[26:4];
  /* ../../HW/src/dp/dp_gen.vhd:1181:94  */
  assign n30721_o = n30719_o == 23'b00000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1182:57  */
  assign n30722_o = d_burstpos_end_r[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1181:17  */
  assign n30724_o = n30721_o ? n30722_o : 4'b1111;
  /* ../../HW/src/dp/dp_gen.vhd:1179:17  */
  assign n30726_o = n30718_o ? 4'b0000 : n30724_o;
  /* ../../HW/src/dp/dp_gen.vhd:1188:55  */
  assign n30727_o = d_bufsize_rr[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:1188:36  */
  assign n30728_o = {2'b0, n30727_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1188:111  */
  assign n30729_o = {1'b0, d_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1188:103  */
  assign n30730_o = n30728_o - n30729_o;
  /* ../../HW/src/dp/dp_gen.vhd:1190:41  */
  assign n30732_o = n30730_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1189:17  */
  assign n30733_o = dst_double_rrr ? n30732_o : n30730_o;
  /* ../../HW/src/dp/dp_gen.vhd:1192:29  */
  assign n30735_o = $signed(n30733_o) <= $signed(25'b0000000000000000000000000);
  /* ../../HW/src/dp/dp_gen.vhd:1194:44  */
  assign n30736_o = {21'b0, d_burstpos_end_rr};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1194:42  */
  assign n30737_o = $unsigned(n30733_o) > $unsigned(n30736_o);
  /* ../../HW/src/dp/dp_gen.vhd:1197:59  */
  assign n30738_o = n30733_o[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1194:17  */
  assign n30739_o = n30737_o ? d_burstpos_end_rr : n30738_o;
  /* ../../HW/src/dp/dp_gen.vhd:1192:17  */
  assign n30741_o = n30735_o ? 4'b0000 : n30739_o;
  /* ../../HW/src/dp/dp_gen.vhd:1201:79  */
  assign n30743_o = d_burst_max_r[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:1201:47  */
  assign n30745_o = {1'b0, n30743_o};
  /* ../../HW/src/dp/dp_gen.vhd:1201:109  */
  assign n30746_o = n30745_o - d_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1202:42  */
  assign n30748_o = dst_vector_r == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1203:106  */
  assign n30749_o = n30746_o[23:1];
  /* ../../HW/src/dp/dp_gen.vhd:1205:45  */
  assign n30752_o = dst_vector_r == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1206:106  */
  assign n30753_o = n30746_o[23:2];
  /* ../../HW/src/dp/dp_gen.vhd:1208:45  */
  assign n30756_o = dst_vector_r == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1209:104  */
  assign n30757_o = n30746_o[23:3];
  assign n30759_o = {3'b000, n30757_o};
  /* ../../HW/src/dp/dp_gen.vhd:1208:17  */
  assign n30760_o = n30756_o ? n30759_o : n30746_o;
  assign n30761_o = {2'b00, n30753_o};
  /* ../../HW/src/dp/dp_gen.vhd:1205:17  */
  assign n30762_o = n30752_o ? n30761_o : n30760_o;
  assign n30763_o = {1'b0, n30749_o};
  /* ../../HW/src/dp/dp_gen.vhd:1202:17  */
  assign n30764_o = n30748_o ? n30763_o : n30762_o;
  /* ../../HW/src/dp/dp_gen.vhd:1214:42  */
  assign n30765_o = d_i0_valid & d_i1_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:57  */
  assign n30766_o = n30765_o & d_i2_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:72  */
  assign n30767_o = n30766_o & d_i3_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:87  */
  assign n30768_o = n30767_o & d_i4_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:102  */
  assign n30769_o = n30768_o & d_burst_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1215:29  */
  assign n30770_o = ~d_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:1217:43  */
  assign n30772_o = dst_is_burst_rr & 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:1218:34  */
  assign n30773_o = d_temp3_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1218:79  */
  assign n30775_o = n30773_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1219:34  */
  assign n30776_o = d_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1219:64  */
  assign n30778_o = n30776_o != 5'b11111;
  /* ../../HW/src/dp/dp_gen.vhd:1218:130  */
  assign n30779_o = n30778_o & n30775_o;
  /* ../../HW/src/dp/dp_gen.vhd:1220:50  */
  assign n30780_o = d_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1218:21  */
  assign n30782_o = n30779_o ? n30780_o : 5'b11110;
  /* ../../HW/src/dp/dp_gen.vhd:1224:39  */
  assign n30783_o = d_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1226:42  */
  assign n30784_o = d_burstremain_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1226:93  */
  assign n30786_o = n30784_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1227:57  */
  assign n30787_o = d_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1227:40  */
  assign n30788_o = $unsigned(n30782_o) > $unsigned(n30787_o);
  /* ../../HW/src/dp/dp_gen.vhd:1226:150  */
  assign n30789_o = n30788_o & n30786_o;
  /* ../../HW/src/dp/dp_gen.vhd:1228:60  */
  assign n30790_o = d_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1228:90  */
  assign n30792_o = n30790_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1230:57  */
  assign n30794_o = n30782_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1226:21  */
  assign n30795_o = n30789_o ? n30792_o : n30794_o;
  /* ../../HW/src/dp/dp_gen.vhd:1224:21  */
  assign n30797_o = n30783_o ? 5'b00000 : n30795_o;
  /* ../../HW/src/dp/dp_gen.vhd:1233:39  */
  assign n30798_o = d_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1233:21  */
  assign n30801_o = n30798_o ? 5'b00000 : 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1217:17  */
  assign n30802_o = n30772_o ? n30797_o : n30801_o;
  /* ../../HW/src/dp/dp_gen.vhd:1215:17  */
  assign n30805_o = n30770_o ? 5'b00000 : n30802_o;
  assign n30828_o = {n30540_o, n30536_o, n30532_o};
  /* ../../HW/src/dp/dp_gen.vhd:915:14  */
  assign n30924_o = n30528_o ? n32871_o : n32892_o;
  /* ../../HW/src/dp/dp_gen.vhd:1252:10  */
  always @*
    n31324_burst_min_v = n32420_q; // (isignal)
  initial
    n31324_burst_min_v = 25'bX;
  /* ../../HW/src/dp/dp_gen.vhd:1256:16  */
  assign n31330_o = ~reset_in;
  /* ../../HW/src/dp/dp_gen.vhd:1333:21  */
  assign n31332_o = ~waitreq;
  /* ../../HW/src/dp/dp_gen.vhd:1333:42  */
  assign n31333_o = instruction_valid_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1333:27  */
  assign n31334_o = n31332_o | n31333_o;
  /* ../../HW/src/dp/dp_gen.vhd:1335:16  */
  assign n31338_o = instruction_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1347:65  */
  assign n31339_o = n29602_o[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1348:71  */
  assign n31340_o = n29602_o[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:1349:69  */
  assign n31341_o = n29602_o[72:48];
  /* ../../HW/src/dp/dp_gen.vhd:1350:69  */
  assign n31342_o = n29602_o[97:73];
  /* ../../HW/src/dp/dp_gen.vhd:1351:65  */
  assign n31343_o = n29602_o[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:1352:71  */
  assign n31344_o = n29602_o[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:1353:69  */
  assign n31345_o = n29602_o[170:146];
  /* ../../HW/src/dp/dp_gen.vhd:1354:69  */
  assign n31346_o = n29602_o[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1355:65  */
  assign n31347_o = n29602_o[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:1356:71  */
  assign n31348_o = n29602_o[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:1357:69  */
  assign n31349_o = n29602_o[268:244];
  /* ../../HW/src/dp/dp_gen.vhd:1358:69  */
  assign n31350_o = n29602_o[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1359:65  */
  assign n31351_o = n29602_o[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:1360:71  */
  assign n31352_o = n29602_o[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:1361:69  */
  assign n31353_o = n29602_o[366:342];
  /* ../../HW/src/dp/dp_gen.vhd:1362:69  */
  assign n31354_o = n29602_o[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1363:65  */
  assign n31355_o = n29602_o[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:1364:71  */
  assign n31356_o = n29602_o[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:1365:69  */
  assign n31357_o = n29602_o[464:440];
  /* ../../HW/src/dp/dp_gen.vhd:1366:69  */
  assign n31358_o = n29602_o[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1367:135  */
  assign n31359_o = n29602_o[514:493];
  /* ../../HW/src/dp/dp_gen.vhd:1369:82  */
  assign n31360_o = n29602_o[490];
  /* ../../HW/src/dp/dp_gen.vhd:1369:99  */
  assign n31361_o = src_vector[0];
  /* ../../HW/src/dp/dp_gen.vhd:1369:86  */
  assign n31362_o = n31360_o | n31361_o;
  /* ../../HW/src/dp/dp_gen.vhd:1369:82  */
  assign n31363_o = n29602_o[491];
  /* ../../HW/src/dp/dp_gen.vhd:1369:99  */
  assign n31364_o = src_vector[1];
  /* ../../HW/src/dp/dp_gen.vhd:1369:86  */
  assign n31365_o = n31363_o | n31364_o;
  /* ../../HW/src/dp/dp_gen.vhd:1369:82  */
  assign n31366_o = n29602_o[492];
  /* ../../HW/src/dp/dp_gen.vhd:1369:99  */
  assign n31367_o = src_vector[2];
  /* ../../HW/src/dp/dp_gen.vhd:1369:86  */
  assign n31368_o = n31366_o | n31367_o;
  /* ../../HW/src/dp/dp_gen.vhd:1371:65  */
  assign n31369_o = n29602_o[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1373:65  */
  assign n31370_o = n29602_o[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:1374:61  */
  assign n31371_o = n29602_o[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:1375:71  */
  assign n31372_o = n29602_o[775:752];
  /* ../../HW/src/dp/dp_gen.vhd:1377:32  */
  assign n31374_o = src_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1378:128  */
  assign n31375_o = n29602_o[648:628];
  /* ../../HW/src/dp/dp_gen.vhd:1380:35  */
  assign n31378_o = src_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1381:130  */
  assign n31379_o = n29602_o[648:627];
  /* ../../HW/src/dp/dp_gen.vhd:1383:35  */
  assign n31382_o = src_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1384:130  */
  assign n31383_o = n29602_o[648:626];
  /* ../../HW/src/dp/dp_gen.vhd:1387:66  */
  assign n31385_o = n29602_o[648:625];
  assign n31386_o = {1'b0, n31383_o};
  /* ../../HW/src/dp/dp_gen.vhd:1383:19  */
  assign n31387_o = n31382_o ? n31386_o : n31385_o;
  assign n31388_o = {2'b00, n31379_o};
  /* ../../HW/src/dp/dp_gen.vhd:1380:19  */
  assign n31389_o = n31378_o ? n31388_o : n31387_o;
  assign n31390_o = {3'b000, n31375_o};
  /* ../../HW/src/dp/dp_gen.vhd:1377:19  */
  assign n31391_o = n31374_o ? n31390_o : n31389_o;
  /* ../../HW/src/dp/dp_gen.vhd:1391:59  */
  assign n31392_o = n29602_o[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1391:69  */
  assign n31394_o = n31392_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1393:59  */
  assign n31395_o = n29602_o[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1390:19  */
  assign n31396_o = source_double_precision ? n31394_o : n31395_o;
  /* ../../HW/src/dp/dp_gen.vhd:1397:44  */
  assign n31397_o = n29602_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1397:55  */
  assign n31399_o = n31397_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1397:19  */
  assign n31402_o = n31399_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1402:32  */
  assign n31404_o = src_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1403:41  */
  assign n31405_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1403:44  */
  assign n31407_o = n31405_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1405:44  */
  assign n31408_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1405:47  */
  assign n31410_o = n31408_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1405:22  */
  assign n31413_o = n31410_o ? 24'b000000000000000001000000 : 24'b000000000000100000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1403:22  */
  assign n31415_o = n31407_o ? 24'b000000000000000000001000 : n31413_o;
  /* ../../HW/src/dp/dp_gen.vhd:1410:35  */
  assign n31417_o = src_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1411:41  */
  assign n31418_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1411:44  */
  assign n31420_o = n31418_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1413:44  */
  assign n31421_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1413:47  */
  assign n31423_o = n31421_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1413:22  */
  assign n31426_o = n31423_o ? 24'b000000000000000000100000 : 24'b000000000000010000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1411:22  */
  assign n31428_o = n31420_o ? 24'b000000000000000000000100 : n31426_o;
  /* ../../HW/src/dp/dp_gen.vhd:1418:35  */
  assign n31430_o = src_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1419:41  */
  assign n31431_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1419:44  */
  assign n31433_o = n31431_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1421:44  */
  assign n31434_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1421:47  */
  assign n31436_o = n31434_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1421:22  */
  assign n31439_o = n31436_o ? 24'b000000000000000000010000 : 24'b000000000000001000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1419:22  */
  assign n31441_o = n31433_o ? 24'b000000000000000000000010 : n31439_o;
  /* ../../HW/src/dp/dp_gen.vhd:1427:62  */
  assign n31442_o = n29602_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1418:19  */
  assign n31443_o = n31430_o ? n31441_o : n31442_o;
  /* ../../HW/src/dp/dp_gen.vhd:1410:19  */
  assign n31444_o = n31417_o ? n31428_o : n31443_o;
  /* ../../HW/src/dp/dp_gen.vhd:1402:19  */
  assign n31445_o = n31404_o ? n31415_o : n31444_o;
  /* ../../HW/src/dp/dp_gen.vhd:1431:60  */
  assign n31447_o = n31445_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1430:19  */
  assign n31448_o = source_double_precision ? n31447_o : n31445_o;
  /* ../../HW/src/dp/dp_gen.vhd:1436:63  */
  assign n31449_o = n29603_o[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1437:69  */
  assign n31450_o = n29603_o[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:1438:67  */
  assign n31451_o = n29603_o[72:48];
  /* ../../HW/src/dp/dp_gen.vhd:1439:63  */
  assign n31452_o = n29603_o[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:1440:69  */
  assign n31453_o = n29603_o[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:1441:67  */
  assign n31454_o = n29603_o[170:146];
  /* ../../HW/src/dp/dp_gen.vhd:1442:63  */
  assign n31455_o = n29603_o[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:1443:69  */
  assign n31456_o = n29603_o[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:1444:67  */
  assign n31457_o = n29603_o[268:244];
  /* ../../HW/src/dp/dp_gen.vhd:1445:63  */
  assign n31458_o = n29603_o[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:1446:69  */
  assign n31459_o = n29603_o[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:1447:67  */
  assign n31460_o = n29603_o[366:342];
  /* ../../HW/src/dp/dp_gen.vhd:1448:63  */
  assign n31461_o = n29603_o[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:1449:69  */
  assign n31462_o = n29603_o[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:1450:67  */
  assign n31463_o = n29603_o[464:440];
  /* ../../HW/src/dp/dp_gen.vhd:1451:59  */
  assign n31464_o = n29603_o[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:1452:63  */
  assign n31465_o = n29603_o[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:1454:56  */
  assign n31466_o = n29603_o[564:540];
  /* ../../HW/src/dp/dp_gen.vhd:1455:65  */
  assign n31467_o = n29603_o[564:540];
  /* ../../HW/src/dp/dp_gen.vhd:1456:66  */
  assign n31468_o = n29603_o[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1457:71  */
  assign n31469_o = n29603_o[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1458:69  */
  assign n31470_o = n29603_o[775:752];
  /* ../../HW/src/dp/dp_gen.vhd:1460:32  */
  assign n31472_o = dst_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1461:126  */
  assign n31473_o = n29603_o[648:628];
  /* ../../HW/src/dp/dp_gen.vhd:1463:35  */
  assign n31476_o = dst_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1464:128  */
  assign n31477_o = n29603_o[648:627];
  /* ../../HW/src/dp/dp_gen.vhd:1466:35  */
  assign n31480_o = dst_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1467:128  */
  assign n31481_o = n29603_o[648:626];
  /* ../../HW/src/dp/dp_gen.vhd:1470:64  */
  assign n31483_o = n29603_o[648:625];
  assign n31484_o = {1'b0, n31481_o};
  /* ../../HW/src/dp/dp_gen.vhd:1466:19  */
  assign n31485_o = n31480_o ? n31484_o : n31483_o;
  assign n31486_o = {2'b00, n31477_o};
  /* ../../HW/src/dp/dp_gen.vhd:1463:19  */
  assign n31487_o = n31476_o ? n31486_o : n31485_o;
  assign n31488_o = {3'b000, n31473_o};
  /* ../../HW/src/dp/dp_gen.vhd:1460:19  */
  assign n31489_o = n31472_o ? n31488_o : n31487_o;
  /* ../../HW/src/dp/dp_gen.vhd:1473:42  */
  assign n31490_o = n29603_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1473:53  */
  assign n31492_o = n31490_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1473:19  */
  assign n31495_o = n31492_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1479:32  */
  assign n31497_o = dst_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1480:41  */
  assign n31498_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1480:44  */
  assign n31500_o = n31498_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1482:44  */
  assign n31502_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1482:47  */
  assign n31504_o = n31502_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1482:22  */
  assign n31507_o = n31504_o ? 24'b000000000000000001000000 : 24'b000000000000100000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1480:22  */
  assign n31508_o = n31500_o ? 24'b000000000000000000001000 : n31507_o;
  /* ../../HW/src/dp/dp_gen.vhd:1487:35  */
  assign n31510_o = dst_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1488:41  */
  assign n31511_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1488:44  */
  assign n31513_o = n31511_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1490:44  */
  assign n31515_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1490:47  */
  assign n31517_o = n31515_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1490:22  */
  assign n31520_o = n31517_o ? 24'b000000000000000000100000 : 24'b000000000000010000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1488:22  */
  assign n31521_o = n31513_o ? 24'b000000000000000000000100 : n31520_o;
  /* ../../HW/src/dp/dp_gen.vhd:1495:35  */
  assign n31523_o = dst_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1496:41  */
  assign n31524_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1496:44  */
  assign n31526_o = n31524_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1498:44  */
  assign n31528_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1498:47  */
  assign n31530_o = n31528_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1498:22  */
  assign n31533_o = n31530_o ? 24'b000000000000000000010000 : 24'b000000000000001000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1496:22  */
  assign n31534_o = n31526_o ? 24'b000000000000000000000010 : n31533_o;
  /* ../../HW/src/dp/dp_gen.vhd:1504:70  */
  assign n31535_o = n29603_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1495:19  */
  assign n31536_o = n31523_o ? n31534_o : n31535_o;
  /* ../../HW/src/dp/dp_gen.vhd:1487:19  */
  assign n31537_o = n31510_o ? n31521_o : n31536_o;
  /* ../../HW/src/dp/dp_gen.vhd:1479:19  */
  assign n31538_o = n31497_o ? n31508_o : n31537_o;
  /* ../../HW/src/dp/dp_gen.vhd:1515:48  */
  assign n31540_o = instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1515:19  */
  assign n31542_o = n31540_o ? 1'b0 : instruction_stream_process_in;
  /* ../../HW/src/dp/dp_gen.vhd:1515:19  */
  assign n31544_o = n31540_o ? instruction_stream_process_in : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1526:50  */
  assign n31546_o = instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1526:102  */
  assign n31548_o = instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1526:72  */
  assign n31549_o = n31548_o & n31546_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:47  */
  assign n31550_o = n29602_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:1527:63  */
  assign n31551_o = ~n31550_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:92  */
  assign n31552_o = n29603_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:1527:108  */
  assign n31553_o = ~n31552_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:68  */
  assign n31554_o = n31553_o & n31551_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:22  */
  assign n31557_o = n31554_o ? 2'b00 : 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1532:78  */
  assign n31558_o = ~dest_double_precision;
  /* ../../HW/src/dp/dp_gen.vhd:1532:53  */
  assign n31559_o = n31558_o & source_double_precision;
  /* ../../HW/src/dp/dp_gen.vhd:1534:48  */
  assign n31560_o = ~source_double_precision;
  /* ../../HW/src/dp/dp_gen.vhd:1534:53  */
  assign n31561_o = dest_double_precision & n31560_o;
  /* ../../HW/src/dp/dp_gen.vhd:1534:19  */
  assign n31564_o = n31561_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1532:19  */
  assign n31566_o = n31559_o ? 2'b01 : n31564_o;
  /* ../../HW/src/dp/dp_gen.vhd:1526:19  */
  assign n31567_o = n31549_o ? n31557_o : n31566_o;
  /* ../../HW/src/dp/dp_gen.vhd:1543:32  */
  assign n31569_o = dst_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1545:105  */
  assign n31571_o = instruction_gen_len_in[23:3];
  /* ../../HW/src/dp/dp_gen.vhd:1545:150  */
  assign n31573_o = n31571_o - 21'b000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1546:35  */
  assign n31575_o = dst_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1548:107  */
  assign n31577_o = instruction_gen_len_in[23:2];
  /* ../../HW/src/dp/dp_gen.vhd:1548:154  */
  assign n31579_o = n31577_o - 22'b0000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1549:35  */
  assign n31581_o = dst_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1551:107  */
  assign n31583_o = instruction_gen_len_in[23:1];
  /* ../../HW/src/dp/dp_gen.vhd:1551:154  */
  assign n31585_o = n31583_o - 23'b00000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1553:58  */
  assign n31587_o = instruction_gen_len_in - 24'b000000000000000000000001;
  assign n31588_o = {1'b0, n31585_o};
  /* ../../HW/src/dp/dp_gen.vhd:1549:19  */
  assign n31589_o = n31581_o ? n31588_o : n31587_o;
  assign n31590_o = {2'b00, n31579_o};
  /* ../../HW/src/dp/dp_gen.vhd:1546:19  */
  assign n31591_o = n31575_o ? n31590_o : n31589_o;
  assign n31592_o = {3'b000, n31573_o};
  /* ../../HW/src/dp/dp_gen.vhd:1543:19  */
  assign n31593_o = n31569_o ? n31592_o : n31591_o;
  /* ../../HW/src/dp/dp_gen.vhd:1557:42  */
  assign n31595_o = n31593_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1557:19  */
  assign n31598_o = n31595_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1572:52  */
  assign n31599_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1573:52  */
  assign n31600_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1572:91  */
  assign n31601_o = {n31599_o, n31600_o};
  /* ../../HW/src/dp/dp_gen.vhd:1574:52  */
  assign n31602_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1573:80  */
  assign n31603_o = {n31601_o, n31602_o};
  /* ../../HW/src/dp/dp_gen.vhd:1575:52  */
  assign n31604_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1574:91  */
  assign n31605_o = {n31603_o, n31604_o};
  /* ../../HW/src/dp/dp_gen.vhd:1576:52  */
  assign n31606_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1575:80  */
  assign n31607_o = {n31605_o, n31606_o};
  /* ../../HW/src/dp/dp_gen.vhd:1577:52  */
  assign n31608_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1576:91  */
  assign n31609_o = {n31607_o, n31608_o};
  /* ../../HW/src/dp/dp_gen.vhd:1578:52  */
  assign n31610_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1577:80  */
  assign n31611_o = {n31609_o, n31610_o};
  /* ../../HW/src/dp/dp_gen.vhd:1579:52  */
  assign n31612_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1578:91  */
  assign n31613_o = {n31611_o, n31612_o};
  /* ../../HW/src/dp/dp_gen.vhd:1581:52  */
  assign n31614_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1582:52  */
  assign n31615_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1581:78  */
  assign n31616_o = {n31614_o, n31615_o};
  /* ../../HW/src/dp/dp_gen.vhd:1583:52  */
  assign n31617_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1582:78  */
  assign n31618_o = {n31616_o, n31617_o};
  /* ../../HW/src/dp/dp_gen.vhd:1584:52  */
  assign n31619_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1583:78  */
  assign n31620_o = {n31618_o, n31619_o};
  /* ../../HW/src/dp/dp_gen.vhd:1585:52  */
  assign n31621_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1584:78  */
  assign n31622_o = {n31620_o, n31621_o};
  /* ../../HW/src/dp/dp_gen.vhd:1586:52  */
  assign n31623_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1585:78  */
  assign n31624_o = {n31622_o, n31623_o};
  /* ../../HW/src/dp/dp_gen.vhd:1587:52  */
  assign n31625_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1586:78  */
  assign n31626_o = {n31624_o, n31625_o};
  /* ../../HW/src/dp/dp_gen.vhd:1588:52  */
  assign n31627_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1587:78  */
  assign n31628_o = {n31626_o, n31627_o};
  /* ../../HW/src/dp/dp_gen.vhd:1571:19  */
  assign n31629_o = source_double_precision ? n31613_o : n31628_o;
  /* ../../HW/src/dp/dp_gen.vhd:1592:44  */
  assign n31630_o = n29602_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1592:55  */
  assign n31632_o = n31630_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1592:19  */
  assign n31635_o = n31632_o ? 1'b1 : 1'b0;
  assign n31636_o = {n31359_o, n31368_o, n31365_o, n31362_o, n31358_o, n31357_o, n31356_o, n31355_o, n31354_o, n31353_o, n31352_o, n31351_o, n31350_o, n31349_o, n31348_o, n31347_o, n31346_o, n31345_o, n31344_o, n31343_o, n31342_o, n31341_o, n31340_o, n31339_o};
  assign n31637_o = {n31445_o, n31391_o, n31371_o, n31396_o};
  assign n31638_o = {n31372_o, n31370_o};
  assign n31646_o = {n31451_o, n31450_o, n31449_o};
  assign n31647_o = {n31454_o, n31453_o, n31452_o};
  assign n31648_o = {n31457_o, n31456_o, n31455_o};
  assign n31649_o = {n31460_o, n31459_o, n31458_o};
  assign n31650_o = {n31463_o, n31462_o, n31461_o};
  assign n31651_o = {n31468_o, n31467_o};
  assign n31652_o = {n31538_o, n31489_o, n31464_o};
  assign n31653_o = {n31470_o, n31465_o};
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n31672_o = instruction_latch_in ? n31466_o : d_burst_max_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n31673_o = instruction_latch_in ? n31593_o : currlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n31684_o = instruction_latch_in ? n31635_o : eof_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n31685_o = instruction_latch_in ? n31598_o : done_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n31703_o = instruction_latch_in ? n31396_o : n31324_burst_min_v;
  /* ../../HW/src/dp/dp_gen.vhd:1614:54  */
  assign n31706_o = n29602_o[97:73];
  /* ../../HW/src/dp/dp_gen.vhd:1615:54  */
  assign n31707_o = n29602_o[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1616:54  */
  assign n31708_o = n29602_o[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1617:54  */
  assign n31709_o = n29602_o[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1618:54  */
  assign n31710_o = n29602_o[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1638:40  */
  assign n31712_o = currlen_new == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1638:16  */
  assign n31715_o = n31712_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1643:34  */
  assign n31716_o = ~s_burstlen_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1647:31  */
  assign n31717_o = ~s_i4_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1652:63  */
  assign n31718_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1654:31  */
  assign n31719_o = ~s_i3_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1661:63  */
  assign n31720_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1662:59  */
  assign n31721_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1664:31  */
  assign n31722_o = ~s_i2_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1673:63  */
  assign n31723_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1674:59  */
  assign n31724_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1675:59  */
  assign n31725_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1677:31  */
  assign n31726_o = ~s_i1_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1689:63  */
  assign n31727_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1690:59  */
  assign n31728_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1691:59  */
  assign n31729_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1692:59  */
  assign n31730_o = s_template_r[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1694:31  */
  assign n31731_o = ~s_i0_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1708:63  */
  assign n31732_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1709:59  */
  assign n31733_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1710:59  */
  assign n31734_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1711:59  */
  assign n31735_o = s_template_r[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1712:59  */
  assign n31736_o = s_template_r[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1715:28  */
  assign n31737_o = ~repeat_r;
  /* ../../HW/src/dp/dp_gen.vhd:1728:63  */
  assign n31738_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1729:59  */
  assign n31739_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1730:59  */
  assign n31740_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1731:59  */
  assign n31741_o = s_template_r[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1732:59  */
  assign n31742_o = s_template_r[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1733:59  */
  assign n31743_o = s_template_r[97:73];
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31745_o = n31731_o ? s_i0_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31747_o = n31731_o ? s_i0_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31748_o = n31731_o ? s_i0_start_new : n31743_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31749_o = n31731_o ? n31736_o : n31742_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31750_o = n31731_o ? n31735_o : n31741_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31751_o = n31731_o ? n31734_o : n31740_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31752_o = n31731_o ? n31733_o : n31739_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31753_o = n31731_o ? n31732_o : n31738_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n31754_o = n31731_o ? eof_r : n31737_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31755_o = n31726_o ? s_i0_r : n31745_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31757_o = n31726_o ? s_i1_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31758_o = n31726_o ? s_i0_count_r : n31747_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31760_o = n31726_o ? s_i1_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31761_o = n31726_o ? s_i0_start_r : n31748_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31762_o = n31726_o ? s_i1_start_new : n31749_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31763_o = n31726_o ? n31730_o : n31750_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31764_o = n31726_o ? n31729_o : n31751_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31765_o = n31726_o ? n31728_o : n31752_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31766_o = n31726_o ? n31727_o : n31753_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n31767_o = n31726_o ? eof_r : n31754_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31768_o = n31722_o ? s_i0_r : n31755_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31769_o = n31722_o ? s_i1_r : n31757_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31771_o = n31722_o ? s_i2_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31772_o = n31722_o ? s_i0_count_r : n31758_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31773_o = n31722_o ? s_i1_count_r : n31760_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31775_o = n31722_o ? s_i2_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31776_o = n31722_o ? s_i0_start_r : n31761_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31777_o = n31722_o ? s_i1_start_r : n31762_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31778_o = n31722_o ? s_i2_start_new : n31763_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31779_o = n31722_o ? n31725_o : n31764_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31780_o = n31722_o ? n31724_o : n31765_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31781_o = n31722_o ? n31723_o : n31766_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n31782_o = n31722_o ? eof_r : n31767_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31783_o = n31719_o ? s_i0_r : n31768_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31784_o = n31719_o ? s_i1_r : n31769_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31785_o = n31719_o ? s_i2_r : n31771_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31787_o = n31719_o ? s_i3_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31788_o = n31719_o ? s_i0_count_r : n31772_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31789_o = n31719_o ? s_i1_count_r : n31773_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31790_o = n31719_o ? s_i2_count_r : n31775_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31792_o = n31719_o ? s_i3_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31793_o = n31719_o ? s_i0_start_r : n31776_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31794_o = n31719_o ? s_i1_start_r : n31777_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31795_o = n31719_o ? s_i2_start_r : n31778_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31796_o = n31719_o ? s_i3_start_new : n31779_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31797_o = n31719_o ? n31721_o : n31780_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31798_o = n31719_o ? n31720_o : n31781_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n31799_o = n31719_o ? eof_r : n31782_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31800_o = n31717_o ? s_i0_r : n31783_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31801_o = n31717_o ? s_i1_r : n31784_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31802_o = n31717_o ? s_i2_r : n31785_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31803_o = n31717_o ? s_i3_r : n31787_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31805_o = n31717_o ? s_i4_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31806_o = n31717_o ? s_i0_count_r : n31788_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31807_o = n31717_o ? s_i1_count_r : n31789_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31808_o = n31717_o ? s_i2_count_r : n31790_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31809_o = n31717_o ? s_i3_count_r : n31792_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31811_o = n31717_o ? s_i4_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31812_o = n31717_o ? s_i0_start_r : n31793_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31813_o = n31717_o ? s_i1_start_r : n31794_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31814_o = n31717_o ? s_i2_start_r : n31795_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31815_o = n31717_o ? s_i3_start_r : n31796_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31816_o = n31717_o ? s_i4_start_new : n31797_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31817_o = n31717_o ? n31718_o : n31798_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n31818_o = n31717_o ? eof_r : n31799_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31819_o = n31716_o ? s_i0_r : n31800_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31820_o = n31716_o ? s_i1_r : n31801_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31821_o = n31716_o ? s_i2_r : n31802_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31822_o = n31716_o ? s_i3_r : n31803_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31823_o = n31716_o ? s_i4_r : n31805_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31824_o = n31716_o ? s_i0_count_r : n31806_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31825_o = n31716_o ? s_i1_count_r : n31807_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31826_o = n31716_o ? s_i2_count_r : n31808_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31827_o = n31716_o ? s_i3_count_r : n31809_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31828_o = n31716_o ? s_i4_count_r : n31811_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31830_o = n31716_o ? s_burstlen_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31832_o = n31716_o ? s_burstpos_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31833_o = n31716_o ? s_i0_start_r : n31812_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31834_o = n31716_o ? s_i1_start_r : n31813_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31835_o = n31716_o ? s_i2_start_r : n31814_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31836_o = n31716_o ? s_i3_start_r : n31815_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31837_o = n31716_o ? s_i4_start_r : n31816_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31838_o = n31716_o ? s_burstpos_start_new : n31817_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n31839_o = n31716_o ? eof_r : n31818_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:34  */
  assign n31840_o = ~d_burstlen_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1738:31  */
  assign n31841_o = ~d_i4_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1743:36  */
  assign n31842_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1743:51  */
  assign n31844_o = n31842_o == 3'b100;
  /* ../../HW/src/dp/dp_gen.vhd:1744:59  */
  assign n31845_o = d_template_r[463:440];
  /* ../../HW/src/dp/dp_gen.vhd:1744:33  */
  assign n31846_o = $unsigned(d_i4_new2) > $unsigned(n31845_o);
  /* ../../HW/src/dp/dp_gen.vhd:1743:55  */
  assign n31847_o = n31846_o & n31844_o;
  /* ../../HW/src/dp/dp_gen.vhd:1745:53  */
  assign n31848_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1747:53  */
  assign n31849_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1743:19  */
  assign n31850_o = n31847_o ? n31848_o : n31849_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:31  */
  assign n31851_o = ~d_i3_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1757:36  */
  assign n31853_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1757:51  */
  assign n31855_o = n31853_o == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1758:59  */
  assign n31856_o = d_template_r[365:342];
  /* ../../HW/src/dp/dp_gen.vhd:1758:33  */
  assign n31857_o = $unsigned(d_i3_new2) > $unsigned(n31856_o);
  /* ../../HW/src/dp/dp_gen.vhd:1757:55  */
  assign n31858_o = n31857_o & n31855_o;
  /* ../../HW/src/dp/dp_gen.vhd:1759:53  */
  assign n31859_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1761:53  */
  assign n31860_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1757:19  */
  assign n31861_o = n31858_o ? n31859_o : n31860_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:31  */
  assign n31862_o = ~d_i2_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1773:36  */
  assign n31864_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1773:51  */
  assign n31866_o = n31864_o == 3'b010;
  /* ../../HW/src/dp/dp_gen.vhd:1774:59  */
  assign n31867_o = d_template_r[267:244];
  /* ../../HW/src/dp/dp_gen.vhd:1774:33  */
  assign n31868_o = $unsigned(d_i2_new2) > $unsigned(n31867_o);
  /* ../../HW/src/dp/dp_gen.vhd:1773:55  */
  assign n31869_o = n31868_o & n31866_o;
  /* ../../HW/src/dp/dp_gen.vhd:1775:53  */
  assign n31870_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1777:53  */
  assign n31871_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1773:19  */
  assign n31872_o = n31869_o ? n31870_o : n31871_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:31  */
  assign n31873_o = ~d_i1_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1791:36  */
  assign n31875_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1791:51  */
  assign n31877_o = n31875_o == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1792:59  */
  assign n31878_o = d_template_r[169:146];
  /* ../../HW/src/dp/dp_gen.vhd:1792:33  */
  assign n31879_o = $unsigned(d_i1_new2) > $unsigned(n31878_o);
  /* ../../HW/src/dp/dp_gen.vhd:1791:55  */
  assign n31880_o = n31879_o & n31877_o;
  /* ../../HW/src/dp/dp_gen.vhd:1793:52  */
  assign n31881_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1795:52  */
  assign n31882_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1791:19  */
  assign n31883_o = n31880_o ? n31881_o : n31882_o;
  /* ../../HW/src/dp/dp_gen.vhd:1797:31  */
  assign n31884_o = ~d_i0_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1811:36  */
  assign n31886_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1811:51  */
  assign n31888_o = n31886_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:1812:59  */
  assign n31889_o = d_template_r[71:48];
  /* ../../HW/src/dp/dp_gen.vhd:1812:33  */
  assign n31890_o = $unsigned(d_i0_new2) > $unsigned(n31889_o);
  /* ../../HW/src/dp/dp_gen.vhd:1811:55  */
  assign n31891_o = n31890_o & n31888_o;
  /* ../../HW/src/dp/dp_gen.vhd:1813:53  */
  assign n31892_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1815:53  */
  assign n31893_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n31894_o = n31900_o ? n31892_o : n31893_o;
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n31897_o = n31884_o ? d_i0_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n31899_o = n31884_o ? d_i0_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n31900_o = n31891_o & n31884_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n31901_o = n31873_o ? d_i0_r : n31897_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n31903_o = n31873_o ? d_i1_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n31904_o = n31873_o ? d_i0_count_r : n31899_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n31906_o = n31873_o ? d_i1_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n31907_o = n31873_o ? n31883_o : n31894_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31908_o = n31862_o ? d_i0_r : n31901_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31909_o = n31862_o ? d_i1_r : n31903_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31911_o = n31862_o ? d_i2_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31912_o = n31862_o ? d_i0_count_r : n31904_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31913_o = n31862_o ? d_i1_count_r : n31906_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31915_o = n31862_o ? d_i2_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n31916_o = n31862_o ? n31872_o : n31907_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31917_o = n31851_o ? d_i0_r : n31908_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31918_o = n31851_o ? d_i1_r : n31909_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31919_o = n31851_o ? d_i2_r : n31911_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31921_o = n31851_o ? d_i3_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31922_o = n31851_o ? d_i0_count_r : n31912_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31923_o = n31851_o ? d_i1_count_r : n31913_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31924_o = n31851_o ? d_i2_count_r : n31915_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31926_o = n31851_o ? d_i3_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n31927_o = n31851_o ? n31861_o : n31916_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31928_o = n31841_o ? d_i0_r : n31917_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31929_o = n31841_o ? d_i1_r : n31918_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31930_o = n31841_o ? d_i2_r : n31919_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31931_o = n31841_o ? d_i3_r : n31921_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31933_o = n31841_o ? d_i4_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31934_o = n31841_o ? d_i0_count_r : n31922_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31935_o = n31841_o ? d_i1_count_r : n31923_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31936_o = n31841_o ? d_i2_count_r : n31924_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31937_o = n31841_o ? d_i3_count_r : n31926_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31939_o = n31841_o ? d_i4_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n31940_o = n31841_o ? n31850_o : n31927_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31941_o = n31840_o ? d_i0_r : n31928_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31942_o = n31840_o ? d_i1_r : n31929_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31943_o = n31840_o ? d_i2_r : n31930_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31944_o = n31840_o ? d_i3_r : n31931_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31945_o = n31840_o ? d_i4_r : n31933_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31946_o = n31840_o ? d_i0_count_r : n31934_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31947_o = n31840_o ? d_i1_count_r : n31935_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31948_o = n31840_o ? d_i2_count_r : n31936_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31949_o = n31840_o ? d_i3_count_r : n31937_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31950_o = n31840_o ? d_i4_count_r : n31939_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31951_o = n31840_o ? d_burst_max_r : n31940_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31953_o = n31840_o ? d_burstlen_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n31955_o = n31840_o ? d_burstpos_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31957_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31959_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31961_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31963_o = reload ? 24'b000000000000000000000000 : n31819_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31965_o = reload ? 24'b000000000000000000000000 : n31820_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31967_o = reload ? 24'b000000000000000000000000 : n31821_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31969_o = reload ? 24'b000000000000000000000000 : n31822_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31971_o = reload ? 24'b000000000000000000000000 : n31823_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31973_o = reload ? 24'b000000000000000000000000 : n31824_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31975_o = reload ? 24'b000000000000000000000000 : n31825_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31977_o = reload ? 24'b000000000000000000000000 : n31826_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31979_o = reload ? 24'b000000000000000000000000 : n31827_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31981_o = reload ? 24'b000000000000000000000000 : n31828_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31983_o = reload ? 24'b000000000000000000000000 : n31830_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31985_o = reload ? 24'b000000000000000000000000 : n31832_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31986_o = reload ? n31706_o : n31833_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31987_o = reload ? n31707_o : n31834_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31988_o = reload ? n31708_o : n31835_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31989_o = reload ? n31709_o : n31836_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31990_o = reload ? n31710_o : n31837_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31991_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31992_o = reload ? n31703_o : n31838_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31994_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31996_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n31998_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32000_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32002_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32004_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32006_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32008_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32010_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32012_o = reload ? 24'b000000000000000000000000 : n31941_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32014_o = reload ? 24'b000000000000000000000000 : n31942_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32016_o = reload ? 24'b000000000000000000000000 : n31943_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32018_o = reload ? 24'b000000000000000000000000 : n31944_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32020_o = reload ? 24'b000000000000000000000000 : n31945_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32022_o = reload ? 24'b000000000000000000000000 : n31946_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32024_o = reload ? 24'b000000000000000000000000 : n31947_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32026_o = reload ? 24'b000000000000000000000000 : n31948_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32028_o = reload ? 24'b000000000000000000000000 : n31949_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32030_o = reload ? 24'b000000000000000000000000 : n31950_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32031_o = reload ? n31672_o : n31951_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32033_o = reload ? 24'b000000000000000000000000 : n31953_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32035_o = reload ? 24'b000000000000000000000000 : n31955_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32036_o = reload ? n31673_o : currlen_new;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32039_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32040_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32041_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32042_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32043_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32044_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32045_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32046_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32047_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32048_o = reload ? n31684_o : n31839_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32049_o = reload ? n31685_o : n31715_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32050_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32051_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32052_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32053_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32054_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32055_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32056_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32057_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32058_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32059_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32060_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32061_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32062_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32063_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32064_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32065_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32066_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32067_o = instruction_valid_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n32069_o = reload ? n31338_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32074_o = n31957_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32076_o = n31959_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32078_o = n31961_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32096_o = n31991_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32099_o = n31994_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32101_o = n31996_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32103_o = n31998_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32105_o = n32000_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32107_o = n32002_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32109_o = n32004_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32111_o = n32006_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32113_o = n32008_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32115_o = n32010_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32131_o = reload & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32132_o = n32039_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32133_o = n32040_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32134_o = n32041_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32135_o = n32042_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32136_o = n32043_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32137_o = n32044_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32138_o = n32045_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32139_o = n32046_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32140_o = n32047_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32143_o = n32050_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32144_o = n32051_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32145_o = n32052_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32146_o = n32053_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32147_o = n32054_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32148_o = n32055_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32149_o = n32056_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32150_o = n32057_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32151_o = n32058_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32152_o = n32059_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32153_o = n32060_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32154_o = n32061_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32155_o = n32062_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32156_o = n32063_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32157_o = n32064_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32158_o = n32065_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32159_o = n32066_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32160_o = n32067_o & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32162_o = n31334_o ? n32069_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n32164_o = reload & n31334_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32417_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32418_o = n32164_o & n32417_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32419_o = n32418_o ? n31703_o : n31324_burst_min_v;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32420_q <= n32419_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32429_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32430_o = n32078_o & n32429_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32431_o = s_template_r[775:728];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32432_o = n32430_o ? n31638_o : n32431_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32433_q <= n32432_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32434_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32435_o = n32076_o & n32434_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32436_o = s_template_r[672:568];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32437_o = n32435_o ? n31637_o : n32436_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32438_q <= n32437_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32439_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32440_o = n32074_o & n32439_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32441_o = s_template_r[514:0];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32442_o = n32440_o ? n31636_o : n32441_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32443_q <= n32442_o;
  assign n32446_o = {n32433_q, 55'bZ, n32438_q, 53'bZ, n32443_q};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32447_o = n31334_o ? n31963_o : s_i0_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32448_q <= 24'b000000000000000000000000;
    else
      n32448_q <= n32447_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32449_o = n31334_o ? n31965_o : s_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32450_q <= 24'b000000000000000000000000;
    else
      n32450_q <= n32449_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32451_o = n31334_o ? n31967_o : s_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32452_q <= 24'b000000000000000000000000;
    else
      n32452_q <= n32451_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32453_o = n31334_o ? n31969_o : s_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32454_q <= 24'b000000000000000000000000;
    else
      n32454_q <= n32453_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32455_o = n31334_o ? n31971_o : s_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32456_q <= 24'b000000000000000000000000;
    else
      n32456_q <= n32455_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32457_o = n31334_o ? n31973_o : s_i0_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32458_q <= 24'b000000000000000000000000;
    else
      n32458_q <= n32457_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32459_o = n31334_o ? n31975_o : s_i1_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32460_q <= 24'b000000000000000000000000;
    else
      n32460_q <= n32459_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32461_o = n31334_o ? n31977_o : s_i2_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32462_q <= 24'b000000000000000000000000;
    else
      n32462_q <= n32461_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32463_o = n31334_o ? n31979_o : s_i3_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32464_q <= 24'b000000000000000000000000;
    else
      n32464_q <= n32463_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32465_o = n31334_o ? n31981_o : s_i4_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32466_q <= 24'b000000000000000000000000;
    else
      n32466_q <= n32465_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32467_o = n31334_o ? n31983_o : s_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32468_q <= 24'b000000000000000000000000;
    else
      n32468_q <= n32467_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32469_o = n31334_o ? n31985_o : s_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32470_q <= 24'b000000000000000000000000;
    else
      n32470_q <= n32469_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32473_o = n30528_o ? n30626_o : s_burstremain_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32474_q <= 24'b111111111111111111111111;
    else
      n32474_q <= n32473_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32475_o = n30528_o ? n30637_o : s_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32476_q <= 1'b1;
    else
      n32476_q <= n32475_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32477_o = n31334_o ? n31986_o : s_i0_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32478_q <= 25'b0000000000000000000000000;
    else
      n32478_q <= n32477_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32479_o = n31334_o ? n31987_o : s_i1_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32480_q <= 25'b0000000000000000000000000;
    else
      n32480_q <= n32479_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32481_o = n31334_o ? n31988_o : s_i2_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32482_q <= 25'b0000000000000000000000000;
    else
      n32482_q <= n32481_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32483_o = n31334_o ? n31989_o : s_i3_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32484_q <= 25'b0000000000000000000000000;
    else
      n32484_q <= n32483_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32485_o = n31334_o ? n31990_o : s_i4_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32486_q <= 25'b0000000000000000000000000;
    else
      n32486_q <= n32485_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32487_o = n32096_o ? n31448_o : s_burstpos_stride_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32488_q <= 24'b000000000000000000000000;
    else
      n32488_q <= n32487_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32489_o = n31334_o ? n31992_o : s_burstpos_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32490_q <= 25'b0000000000000000000000000;
    else
      n32490_q <= n32489_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32491_o = n30528_o ? n30690_o : s_burstpos_start_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32492_q <= 4'b0000;
    else
      n32492_q <= n32491_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32493_o = n30528_o ? s_burstpos_start_rr : s_burstpos_start_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32494_q <= 4'b0000;
    else
      n32494_q <= n32493_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32495_o = n30528_o ? s_burstpos_start_rrr : s_burstpos_start_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32496_q <= 4'b0000;
    else
      n32496_q <= n32495_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32497_o = n30528_o ? n30579_o : s_burstpos_end_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32498_q <= 27'b000000000000000000000000000;
    else
      n32498_q <= n32497_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32499_o = n30528_o ? n30588_o : s_burstpos_end_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32500_q <= 4'b0000;
    else
      n32500_q <= n32499_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32501_o = n30528_o ? n30603_o : s_burstpos_end_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32502_q <= 4'b0000;
    else
      n32502_q <= n32501_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32503_o = n30528_o ? n30717_o : d_burstpos_end_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32504_q <= 27'b000000000000000000000000000;
    else
      n32504_q <= n32503_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32505_o = n30528_o ? n30726_o : d_burstpos_end_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32506_q <= 4'b0000;
    else
      n32506_q <= n32505_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32507_o = n30528_o ? n30741_o : d_burstpos_end_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32508_q <= 4'b0000;
    else
      n32508_q <= n32507_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32509_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32510_o = n32115_o & n32509_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32511_o = d_template_r[775:728];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32512_o = n32510_o ? n31653_o : n32511_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32513_q <= n32512_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32514_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32515_o = n32113_o & n32514_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32516_o = d_template_r[672:593];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32517_o = n32515_o ? n31652_o : n32516_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32518_q <= n32517_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32519_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32520_o = n32111_o & n32519_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32521_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32522_o = n32520_o ? n31469_o : n32521_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32523_q <= n32522_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32524_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32525_o = n32109_o & n32524_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32526_o = d_template_r[539:490];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32527_o = n32525_o ? n31651_o : n32526_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32528_q <= n32527_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32529_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32530_o = n32107_o & n32529_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32531_o = d_template_r[464:392];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32532_o = n32530_o ? n31650_o : n32531_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32533_q <= n32532_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32534_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32535_o = n32105_o & n32534_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32536_o = d_template_r[366:294];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32537_o = n32535_o ? n31649_o : n32536_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32538_q <= n32537_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32539_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32540_o = n32103_o & n32539_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32541_o = d_template_r[268:196];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32542_o = n32540_o ? n31648_o : n32541_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32543_q <= n32542_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32544_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32545_o = n32101_o & n32544_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32546_o = d_template_r[170:98];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32547_o = n32545_o ? n31647_o : n32546_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32548_q <= n32547_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32549_o = ~n31330_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n32550_o = n32099_o & n32549_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32551_o = d_template_r[72:0];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32552_o = n32550_o ? n31646_o : n32551_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n32553_q <= n32552_o;
  assign n32562_o = {n32513_q, 55'bZ, n32518_q, 25'bZ, n32523_q, 25'bZ, n32528_q, 25'bZ, n32533_q, 25'bZ, n32538_q, 25'bZ, n32543_q, 25'bZ, n32548_q, 25'bZ, n32553_q};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32563_o = n31334_o ? n32012_o : d_i0_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32564_q <= 24'b000000000000000000000000;
    else
      n32564_q <= n32563_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32565_o = n31334_o ? n32014_o : d_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32566_q <= 24'b000000000000000000000000;
    else
      n32566_q <= n32565_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32567_o = n31334_o ? n32016_o : d_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32568_q <= 24'b000000000000000000000000;
    else
      n32568_q <= n32567_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32569_o = n31334_o ? n32018_o : d_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32570_q <= 24'b000000000000000000000000;
    else
      n32570_q <= n32569_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32571_o = n31334_o ? n32020_o : d_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32572_q <= 24'b000000000000000000000000;
    else
      n32572_q <= n32571_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32573_o = n31334_o ? n32022_o : d_i0_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32574_q <= 24'b000000000000000000000000;
    else
      n32574_q <= n32573_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32575_o = n31334_o ? n32024_o : d_i1_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32576_q <= 24'b000000000000000000000000;
    else
      n32576_q <= n32575_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32577_o = n31334_o ? n32026_o : d_i2_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32578_q <= 24'b000000000000000000000000;
    else
      n32578_q <= n32577_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32579_o = n31334_o ? n32028_o : d_i3_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32580_q <= 24'b000000000000000000000000;
    else
      n32580_q <= n32579_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32581_o = n31334_o ? n32030_o : d_i4_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32582_q <= 24'b000000000000000000000000;
    else
      n32582_q <= n32581_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32583_o = n31334_o ? n32031_o : d_burst_max_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32584_q <= 25'b0000000000000000000000000;
    else
      n32584_q <= n32583_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32585_o = n31334_o ? n32033_o : d_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32586_q <= 24'b000000000000000000000000;
    else
      n32586_q <= n32585_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32587_o = n31334_o ? n32035_o : d_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32588_q <= 24'b000000000000000000000000;
    else
      n32588_q <= n32587_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32591_o = n30528_o ? n30764_o : d_burstremain_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32592_q <= 24'b111111111111111111111111;
    else
      n32592_q <= n32591_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32593_o = n30528_o ? n30769_o : d_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32594_q <= 1'b1;
    else
      n32594_q <= n32593_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32595_o = n31334_o ? n32036_o : currlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32596_q <= 24'b000000000000000000000000;
    else
      n32596_q <= n32595_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32599_o = n32131_o ? instruction_valid_in : running_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32600_q <= 1'b0;
    else
      n32600_q <= n32599_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32601_o = n30528_o ? running_r : running_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32602_q <= 1'b0;
    else
      n32602_q <= n32601_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32603_o = n30528_o ? running_rr : running_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32604_q <= 1'b0;
    else
      n32604_q <= n32603_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32605_o = n30528_o ? running_rrr : running_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32606_q <= 1'b0;
    else
      n32606_q <= n32605_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32607_o = n30528_o ? n30828_o : gen_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32608_q <= 3'b000;
    else
      n32608_q <= n32607_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32609_o = n32132_o ? instruction_bus_id_dest_in : dp_dst_bus_id_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32610_q <= 2'b00;
    else
      n32610_q <= n32609_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32611_o = n30528_o ? dp_dst_bus_id_r : dp_dst_bus_id_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32612_q <= 2'b00;
    else
      n32612_q <= n32611_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32613_o = n30528_o ? dp_dst_bus_id_rr : dp_dst_bus_id_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32614_q <= 2'b00;
    else
      n32614_q <= n32613_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32615_o = n30528_o ? dp_dst_bus_id_rrr : dp_dst_bus_id_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32616_q <= 2'b00;
    else
      n32616_q <= n32615_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32617_o = n32133_o ? instruction_bus_id_source_in : dp_src_bus_id_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32618_q <= 2'b00;
    else
      n32618_q <= n32617_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32619_o = n30528_o ? dp_src_bus_id_r : dp_src_bus_id_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32620_q <= 2'b00;
    else
      n32620_q <= n32619_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32621_o = n30528_o ? dp_src_bus_id_rr : dp_src_bus_id_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32622_q <= 2'b00;
    else
      n32622_q <= n32621_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32623_o = n30528_o ? dp_src_bus_id_rrr : dp_src_bus_id_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32624_q <= 2'b00;
    else
      n32624_q <= n32623_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32625_o = n32134_o ? instruction_data_type_dest_in : dp_dst_data_type_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32626_q <= 2'b00;
    else
      n32626_q <= n32625_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32627_o = n30528_o ? dp_dst_data_type_r : dp_dst_data_type_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32628_q <= 2'b00;
    else
      n32628_q <= n32627_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32629_o = n30528_o ? dp_dst_data_type_rr : dp_dst_data_type_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32630_q <= 2'b00;
    else
      n32630_q <= n32629_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32631_o = n30528_o ? dp_dst_data_type_rrr : dp_dst_data_type_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32632_q <= 2'b00;
    else
      n32632_q <= n32631_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32633_o = n32135_o ? instruction_data_type_source_in : dp_src_data_type_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32634_q <= 2'b00;
    else
      n32634_q <= n32633_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32635_o = n30528_o ? dp_src_data_type_r : dp_src_data_type_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32636_q <= 2'b00;
    else
      n32636_q <= n32635_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32637_o = n30528_o ? dp_src_data_type_rr : dp_src_data_type_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32638_q <= 2'b00;
    else
      n32638_q <= n32637_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32639_o = n30528_o ? dp_src_data_type_rrr : dp_src_data_type_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32640_q <= 2'b00;
    else
      n32640_q <= n32639_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32641_o = n32136_o ? instruction_data_model_source_in : dp_src_data_model_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32642_q <= 2'b00;
    else
      n32642_q <= n32641_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32643_o = n30528_o ? dp_src_data_model_r : dp_src_data_model_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32644_q <= 2'b00;
    else
      n32644_q <= n32643_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32645_o = n30528_o ? dp_src_data_model_rr : dp_src_data_model_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32646_q <= 2'b00;
    else
      n32646_q <= n32645_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32647_o = n30528_o ? dp_src_data_model_rrr : dp_src_data_model_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32648_q <= 2'b00;
    else
      n32648_q <= n32647_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32649_o = n32137_o ? instruction_data_model_dest_in : dp_dst_data_model_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32650_q <= 2'b00;
    else
      n32650_q <= n32649_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32651_o = n30528_o ? dp_dst_data_model_r : dp_dst_data_model_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32652_q <= 2'b00;
    else
      n32652_q <= n32651_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32653_o = n30528_o ? dp_dst_data_model_rr : dp_dst_data_model_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32654_q <= 2'b00;
    else
      n32654_q <= n32653_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32655_o = n30528_o ? dp_dst_data_model_rrr : dp_dst_data_model_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32656_q <= 2'b00;
    else
      n32656_q <= n32655_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32657_o = n32138_o ? instruction_thread_in : dp_thread_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32658_q <= 1'b0;
    else
      n32658_q <= n32657_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32659_o = n30528_o ? dp_thread_r : dp_thread_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32660_q <= 1'b0;
    else
      n32660_q <= n32659_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32661_o = n30528_o ? dp_thread_rr : dp_thread_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32662_q <= 1'b0;
    else
      n32662_q <= n32661_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32663_o = n30528_o ? dp_thread_rrr : dp_thread_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32664_q <= 1'b0;
    else
      n32664_q <= n32663_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32665_o = n32139_o ? instruction_mcast_in : dp_mcast_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32666_q <= 6'b111111;
    else
      n32666_q <= n32665_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32667_o = n30528_o ? dp_mcast_r : dp_mcast_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32668_q <= 6'b111111;
    else
      n32668_q <= n32667_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32669_o = n30528_o ? dp_mcast_rr : dp_mcast_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32670_q <= 6'b111111;
    else
      n32670_q <= n32669_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32671_o = n30528_o ? dp_mcast_rrr : dp_mcast_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32672_q <= 6'b111111;
    else
      n32672_q <= n32671_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32673_o = n32140_o ? n31629_o : data_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32674_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n32674_q <= n32673_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32675_o = n30528_o ? data_r : data_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32676_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n32676_q <= n32675_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32677_o = n30528_o ? data_rr : data_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32678_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n32678_q <= n32677_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32679_o = n30528_o ? data_rrr : data_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32680_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n32680_q <= n32679_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32681_o = n30528_o ? n30546_o : s_bufsize_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32682_q <= 24'b000000000000000000000000;
    else
      n32682_q <= n32681_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32683_o = n30528_o ? s_bufsize_r : s_bufsize_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32684_q <= 24'b000000000000000000000000;
    else
      n32684_q <= n32683_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32685_o = n30528_o ? n30545_o : s_temp1_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32686_q <= 24'b000000000000000000000000;
    else
      n32686_q <= n32685_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32687_o = n30528_o ? n30547_o : s_temp2_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32688_q <= 32'b00000000000000000000000000000000;
    else
      n32688_q <= n32687_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32689_o = n30528_o ? n30549_o : s_temp3_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32690_q <= 24'b000000000000000000000000;
    else
      n32690_q <= n32689_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32691_o = n30528_o ? n30551_o : s_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32692_q <= 24'b000000000000000000000000;
    else
      n32692_q <= n32691_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32693_o = n30528_o ? n30552_o : s_temp5_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32694_q <= 24'b000000000000000000000000;
    else
      n32694_q <= n32693_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32695_o = n30528_o ? s_temp2_r : s_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32696_q <= 32'b00000000000000000000000000000000;
    else
      n32696_q <= n32695_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32697_o = n30528_o ? n30557_o : s_gen_addr_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32698_q <= 32'b00000000000000000000000000000000;
    else
      n32698_q <= n32697_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32699_o = n30528_o ? n30673_o : s_gen_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32700_q <= 5'b00000;
    else
      n32700_q <= n32699_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32701_o = n30528_o ? n30565_o : s_gen_burstlen_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32702_q <= 5'b00000;
    else
      n32702_q <= n32701_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32703_o = n30528_o ? n30570_o : s_gen_burstlen_progress_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32704_q <= 1'b0;
    else
      n32704_q <= n32703_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32705_o = n30528_o ? n30695_o : d_bufsize_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32706_q <= 24'b000000000000000000000000;
    else
      n32706_q <= n32705_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32707_o = n30528_o ? d_bufsize_r : d_bufsize_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32708_q <= 24'b000000000000000000000000;
    else
      n32708_q <= n32707_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32709_o = n30528_o ? n30697_o : d_temp1_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32710_q <= 24'b000000000000000000000000;
    else
      n32710_q <= n32709_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32711_o = n30528_o ? n30698_o : d_temp2_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32712_q <= 32'b00000000000000000000000000000000;
    else
      n32712_q <= n32711_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32713_o = n30528_o ? n30700_o : d_temp3_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32714_q <= 24'b000000000000000000000000;
    else
      n32714_q <= n32713_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32715_o = n30528_o ? n30702_o : d_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32716_q <= 24'b000000000000000000000000;
    else
      n32716_q <= n32715_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32717_o = n30528_o ? n30703_o : d_temp5_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32718_q <= 24'b000000000000000000000000;
    else
      n32718_q <= n32717_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32719_o = n30528_o ? d_temp2_r : d_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32720_q <= 32'b00000000000000000000000000000000;
    else
      n32720_q <= n32719_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32721_o = n30528_o ? n30708_o : d_gen_addr_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32722_q <= 32'b00000000000000000000000000000000;
    else
      n32722_q <= n32721_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32723_o = n30528_o ? n30805_o : d_gen_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32724_q <= 5'b00000;
    else
      n32724_q <= n32723_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32725_o = n30528_o ? d_gen_burstlen_r : d_gen_burstlen_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32726_q <= 5'b00000;
    else
      n32726_q <= n32725_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32727_o = n31334_o ? n32048_o : eof_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32728_q <= 1'b0;
    else
      n32728_q <= n32727_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32729_o = n30528_o ? eof_r : eof_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32730_q <= 1'b0;
    else
      n32730_q <= n32729_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32731_o = n30528_o ? eof_rr : eof_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32732_q <= 1'b0;
    else
      n32732_q <= n32731_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32733_o = n30528_o ? eof_rrr : eof_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32734_q <= 1'b0;
    else
      n32734_q <= n32733_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32735_o = n31334_o ? n32049_o : done_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32736_q <= 1'b1;
    else
      n32736_q <= n32735_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32737_o = n32143_o ? instruction_repeat_in : repeat_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32738_q <= 1'b0;
    else
      n32738_q <= n32737_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32739_o = n32144_o ? n31567_o : data_flow_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32740_q <= 2'b00;
    else
      n32740_q <= n32739_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32741_o = n30528_o ? data_flow_r : data_flow_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32742_q <= 2'b00;
    else
      n32742_q <= n32741_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32743_o = n30528_o ? data_flow_rr : data_flow_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32744_q <= 2'b00;
    else
      n32744_q <= n32743_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32745_o = n30528_o ? data_flow_rrr : data_flow_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32746_q <= 2'b00;
    else
      n32746_q <= n32745_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32747_o = n32145_o ? n31542_o : stream_src_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32748_q <= 1'b0;
    else
      n32748_q <= n32747_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32749_o = n30528_o ? stream_src_r : stream_src_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32750_q <= 1'b0;
    else
      n32750_q <= n32749_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32751_o = n30528_o ? stream_src_rr : stream_src_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32752_q <= 1'b0;
    else
      n32752_q <= n32751_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32753_o = n30528_o ? stream_src_rrr : stream_src_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32754_q <= 1'b0;
    else
      n32754_q <= n32753_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32755_o = n32146_o ? n31544_o : stream_dest_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32756_q <= 1'b0;
    else
      n32756_q <= n32755_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32757_o = n30528_o ? stream_dest_r : stream_dest_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32758_q <= 1'b0;
    else
      n32758_q <= n32757_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32759_o = n30528_o ? stream_dest_rr : stream_dest_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32760_q <= 1'b0;
    else
      n32760_q <= n32759_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32761_o = n30528_o ? stream_dest_rrr : stream_dest_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32762_q <= 1'b0;
    else
      n32762_q <= n32761_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32763_o = n32147_o ? instruction_vm_in : vm_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32764_q <= 1'b0;
    else
      n32764_q <= n32763_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32765_o = n30528_o ? vm_r : vm_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32766_q <= 1'b0;
    else
      n32766_q <= n32765_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32767_o = n30528_o ? vm_rr : vm_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32768_q <= 1'b0;
    else
      n32768_q <= n32767_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32769_o = n30528_o ? vm_rrr : vm_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32770_q <= 1'b0;
    else
      n32770_q <= n32769_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32771_o = n32148_o ? instruction_stream_process_id_in : stream_id_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32772_q <= 2'b00;
    else
      n32772_q <= n32771_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32773_o = n30528_o ? stream_id_r : stream_id_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32774_q <= 2'b00;
    else
      n32774_q <= n32773_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32775_o = n30528_o ? stream_id_rr : stream_id_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32776_q <= 2'b00;
    else
      n32776_q <= n32775_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32777_o = n30528_o ? stream_id_rrr : stream_id_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32778_q <= 2'b00;
    else
      n32778_q <= n32777_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32779_o = n32149_o ? source_double_precision : src_double_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32780_q <= 1'b0;
    else
      n32780_q <= n32779_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32781_o = n30528_o ? src_double_r : src_double_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32782_q <= 1'b0;
    else
      n32782_q <= n32781_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32783_o = n30528_o ? src_double_rr : src_double_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32784_q <= 1'b0;
    else
      n32784_q <= n32783_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32787_o = n32150_o ? dest_double_precision : dst_double_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32788_q <= 1'b0;
    else
      n32788_q <= n32787_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32789_o = n30528_o ? dst_double_r : dst_double_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32790_q <= 1'b0;
    else
      n32790_q <= n32789_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32791_o = n30528_o ? dst_double_rr : dst_double_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32792_q <= 1'b0;
    else
      n32792_q <= n32791_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32795_o = n32151_o ? src_vector : src_vector_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32796_q <= 3'b000;
    else
      n32796_q <= n32795_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32797_o = n30528_o ? src_vector_r : src_vector_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32798_q <= 3'b000;
    else
      n32798_q <= n32797_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32799_o = n30528_o ? src_vector_rr : src_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32800_q <= 3'b000;
    else
      n32800_q <= n32799_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32801_o = n30528_o ? n30678_o : src_vector_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32802_q <= 3'b000;
    else
      n32802_q <= n32801_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32803_o = n32152_o ? dst_vector : dst_vector_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32804_q <= 3'b000;
    else
      n32804_q <= n32803_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32805_o = n30528_o ? dst_vector_r : dst_vector_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32806_q <= 3'b000;
    else
      n32806_q <= n32805_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32807_o = n30528_o ? dst_vector_rr : dst_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32808_q <= 3'b000;
    else
      n32808_q <= n32807_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32809_o = n30528_o ? n30694_o : dst_vector_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32810_q <= 3'b000;
    else
      n32810_q <= n32809_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32811_o = n32153_o ? instruction_source_addr_mode_in : src_addr_mode_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32812_q <= 1'b0;
    else
      n32812_q <= n32811_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32813_o = n30528_o ? src_addr_mode_r : src_addr_mode_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32814_q <= 1'b0;
    else
      n32814_q <= n32813_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32815_o = n30528_o ? src_addr_mode_rr : src_addr_mode_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32816_q <= 1'b0;
    else
      n32816_q <= n32815_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32817_o = n30528_o ? src_addr_mode_rrr : src_addr_mode_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32818_q <= 1'b0;
    else
      n32818_q <= n32817_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32819_o = n32154_o ? instruction_dest_addr_mode_in : dst_addr_mode_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32820_q <= 1'b0;
    else
      n32820_q <= n32819_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32821_o = n30528_o ? dst_addr_mode_r : dst_addr_mode_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32822_q <= 1'b0;
    else
      n32822_q <= n32821_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32823_o = n30528_o ? dst_addr_mode_rr : dst_addr_mode_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32824_q <= 1'b0;
    else
      n32824_q <= n32823_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32825_o = n30528_o ? dst_addr_mode_rrr : dst_addr_mode_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32826_q <= 1'b0;
    else
      n32826_q <= n32825_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32827_o = n32155_o ? src_scatter : src_scatter_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32828_q <= 2'b00;
    else
      n32828_q <= n32827_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32829_o = n30528_o ? src_scatter_r : src_scatter_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32830_q <= 2'b00;
    else
      n32830_q <= n32829_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32831_o = n30528_o ? src_scatter_rr : src_scatter_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32832_q <= 2'b00;
    else
      n32832_q <= n32831_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32833_o = n30528_o ? src_scatter_rrr : src_scatter_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32834_q <= 2'b00;
    else
      n32834_q <= n32833_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32835_o = n32156_o ? dst_scatter : dst_scatter_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32836_q <= 2'b00;
    else
      n32836_q <= n32835_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32837_o = n30528_o ? dst_scatter_r : dst_scatter_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32838_q <= 2'b00;
    else
      n32838_q <= n32837_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32839_o = n30528_o ? dst_scatter_rr : dst_scatter_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32840_q <= 2'b00;
    else
      n32840_q <= n32839_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32841_o = n30528_o ? dst_scatter_rrr : dst_scatter_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32842_q <= 2'b00;
    else
      n32842_q <= n32841_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32843_o = n32157_o ? n31402_o : src_is_burst_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32844_q <= 1'b0;
    else
      n32844_q <= n32843_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32845_o = n30528_o ? src_is_burst_r : src_is_burst_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32846_q <= 1'b0;
    else
      n32846_q <= n32845_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32847_o = n32158_o ? n31495_o : dst_is_burst_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32848_q <= 1'b0;
    else
      n32848_q <= n32847_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n32849_o = n30528_o ? dst_is_burst_r : dst_is_burst_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32850_q <= 1'b0;
    else
      n32850_q <= n32849_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n29686_o)
    if (n29686_o)
      n32852_q <= 3'b000;
    else
      n32852_q <= n30147_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n29686_o)
    if (n29686_o)
      n32853_q <= 3'b000;
    else
      n32853_q <= n30149_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n29686_o)
    if (n29686_o)
      n32854_q <= 6'b000000;
    else
      n32854_q <= n30151_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n29686_o)
    if (n29686_o)
      n32855_q <= 6'b000000;
    else
      n32855_q <= n30153_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32856_o = n32159_o ? n31369_o : s_burst_actual_max_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32857_q <= 25'b0000000000000000000000000;
    else
      n32857_q <= n32856_o;
  /* ../../HW/src/dp/dp_gen.vhd:1256:4  */
  assign n32858_o = {14'b00000000000000, dest_double_precision, dst_scatter, dst_vector, instruction_bus_id_dest_in, source_double_precision, src_scatter, src_vector, instruction_bus_id_source_in, 2'b01};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n32859_o = n32160_o ? log : log_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32860_q <= 32'b00000000000000000000000000000000;
    else
      n32860_q <= n32859_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n31330_o)
    if (n31330_o)
      n32861_q <= 1'b0;
    else
      n32861_q <= n32162_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n30526_o)
    if (n30526_o)
      n32864_q <= 1'b0;
    else
      n32864_q <= n30924_o;
  /* ../../HW/src/dp/dp_gen.vhd:121:16  */
  assign n32865_o = wr_full_in[0];
  /* ../../HW/src/dp/dp_gen.vhd:120:16  */
  assign n32866_o = wr_full_in[1];
  /* ../../HW/src/dp/dp_gen.vhd:116:16  */
  assign n32867_o = wr_full_in[2];
  /* ../../HW/src/dp/dp_gen.vhd:115:16  */
  assign n32868_o = dp_dst_bus_id_rrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:926:46  */
  assign n32869_o = n32868_o ? n32866_o : n32865_o;
  /* ../../HW/src/dp/dp_gen.vhd:113:16  */
  assign n32870_o = dp_dst_bus_id_rrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:926:46  */
  assign n32871_o = n32870_o ? n32867_o : n32869_o;
  /* ../../HW/src/dp/dp_gen.vhd:926:46  */
  assign n32872_o = wr_maxburstlen_in[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:926:47  */
  assign n32873_o = wr_maxburstlen_in[9:5];
  /* ../../HW/src/dp/dp_gen.vhd:111:16  */
  assign n32874_o = wr_maxburstlen_in[14:10];
  /* ../../HW/src/dp/dp_gen.vhd:110:16  */
  assign n32875_o = dp_dst_bus_id_rrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:985:56  */
  assign n32876_o = n32875_o ? n32873_o : n32872_o;
  /* ../../HW/src/dp/dp_gen.vhd:108:16  */
  assign n32877_o = dp_dst_bus_id_rrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:985:56  */
  assign n32878_o = n32877_o ? n32874_o : n32876_o;
  /* ../../HW/src/dp/dp_gen.vhd:985:56  */
  assign n32879_o = wr_maxburstlen_in[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:985:57  */
  assign n32880_o = wr_maxburstlen_in[9:5];
  /* ../../HW/src/dp/dp_gen.vhd:106:16  */
  assign n32881_o = wr_maxburstlen_in[14:10];
  /* ../../HW/src/dp/dp_gen.vhd:105:16  */
  assign n32882_o = dp_dst_bus_id_rrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:986:54  */
  assign n32883_o = n32882_o ? n32880_o : n32879_o;
  /* ../../HW/src/dp/dp_gen.vhd:103:16  */
  assign n32884_o = dp_dst_bus_id_rrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:986:54  */
  assign n32885_o = n32884_o ? n32881_o : n32883_o;
  /* ../../HW/src/dp/dp_gen.vhd:986:54  */
  assign n32886_o = wr_full_in[0];
  /* ../../HW/src/dp/dp_gen.vhd:986:55  */
  assign n32887_o = wr_full_in[1];
  /* ../../HW/src/dp/dp_gen.vhd:101:16  */
  assign n32888_o = wr_full_in[2];
  /* ../../HW/src/dp/dp_gen.vhd:100:16  */
  assign n32889_o = dp_dst_bus_id_rrrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:1240:46  */
  assign n32890_o = n32889_o ? n32887_o : n32886_o;
  /* ../../HW/src/dp/dp_gen.vhd:98:16  */
  assign n32891_o = dp_dst_bus_id_rrrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:1240:46  */
  assign n32892_o = n32891_o ? n32888_o : n32890_o;
endmodule

module dp_gen_3_0_5b55ec37559bb110228a6591713076b7fa2ce5e8
  (input  clock_in,
   input  reset_in,
   input  instruction_valid_in,
   input  instruction_latch_in,
   input  [23:0] instruction_source_in_stride0,
   input  [23:0] instruction_source_in_stride0_count,
   input  [24:0] instruction_source_in_stride0_max,
   input  [24:0] instruction_source_in_stride0_min,
   input  [23:0] instruction_source_in_stride1,
   input  [23:0] instruction_source_in_stride1_count,
   input  [24:0] instruction_source_in_stride1_max,
   input  [24:0] instruction_source_in_stride1_min,
   input  [23:0] instruction_source_in_stride2,
   input  [23:0] instruction_source_in_stride2_count,
   input  [24:0] instruction_source_in_stride2_max,
   input  [24:0] instruction_source_in_stride2_min,
   input  [23:0] instruction_source_in_stride3,
   input  [23:0] instruction_source_in_stride3_count,
   input  [24:0] instruction_source_in_stride3_max,
   input  [24:0] instruction_source_in_stride3_min,
   input  [23:0] instruction_source_in_stride4,
   input  [23:0] instruction_source_in_stride4_count,
   input  [24:0] instruction_source_in_stride4_max,
   input  [24:0] instruction_source_in_stride4_min,
   input  [24:0] instruction_source_in_burst_max,
   input  [24:0] instruction_source_in_burst_max2,
   input  [24:0] instruction_source_in_burst_max_init,
   input  [2:0] instruction_source_in_burst_max_index,
   input  [24:0] instruction_source_in_burst_min,
   input  [31:0] instruction_source_in_bar,
   input  [23:0] instruction_source_in_count,
   input  [23:0] instruction_source_in_burststride,
   input  instruction_source_in_double_precision,
   input  [1:0] instruction_source_in_data_model,
   input  instruction_source_in_scatter,
   input  [23:0] instruction_source_in_totalcount,
   input  [5:0] instruction_source_in_mcast,
   input  [15:0] instruction_source_in_data,
   input  instruction_source_in_repeat,
   input  [1:0] instruction_source_in_datatype,
   input  [1:0] instruction_source_in_bus_id,
   input  [23:0] instruction_source_in_bufsize,
   input  [23:0] instruction_source_in_burst_max_len,
   input  [23:0] instruction_dest_in_stride0,
   input  [23:0] instruction_dest_in_stride0_count,
   input  [24:0] instruction_dest_in_stride0_max,
   input  [24:0] instruction_dest_in_stride0_min,
   input  [23:0] instruction_dest_in_stride1,
   input  [23:0] instruction_dest_in_stride1_count,
   input  [24:0] instruction_dest_in_stride1_max,
   input  [24:0] instruction_dest_in_stride1_min,
   input  [23:0] instruction_dest_in_stride2,
   input  [23:0] instruction_dest_in_stride2_count,
   input  [24:0] instruction_dest_in_stride2_max,
   input  [24:0] instruction_dest_in_stride2_min,
   input  [23:0] instruction_dest_in_stride3,
   input  [23:0] instruction_dest_in_stride3_count,
   input  [24:0] instruction_dest_in_stride3_max,
   input  [24:0] instruction_dest_in_stride3_min,
   input  [23:0] instruction_dest_in_stride4,
   input  [23:0] instruction_dest_in_stride4_count,
   input  [24:0] instruction_dest_in_stride4_max,
   input  [24:0] instruction_dest_in_stride4_min,
   input  [24:0] instruction_dest_in_burst_max,
   input  [24:0] instruction_dest_in_burst_max2,
   input  [24:0] instruction_dest_in_burst_max_init,
   input  [2:0] instruction_dest_in_burst_max_index,
   input  [24:0] instruction_dest_in_burst_min,
   input  [31:0] instruction_dest_in_bar,
   input  [23:0] instruction_dest_in_count,
   input  [23:0] instruction_dest_in_burststride,
   input  instruction_dest_in_double_precision,
   input  [1:0] instruction_dest_in_data_model,
   input  instruction_dest_in_scatter,
   input  [23:0] instruction_dest_in_totalcount,
   input  [5:0] instruction_dest_in_mcast,
   input  [15:0] instruction_dest_in_data,
   input  instruction_dest_in_repeat,
   input  [1:0] instruction_dest_in_datatype,
   input  [1:0] instruction_dest_in_bus_id,
   input  [23:0] instruction_dest_in_bufsize,
   input  [23:0] instruction_dest_in_burst_max_len,
   input  instruction_stream_process_in,
   input  [1:0] instruction_stream_process_id_in,
   input  instruction_vm_in,
   input  [23:0] pre_instruction_source_in_stride0,
   input  [23:0] pre_instruction_source_in_stride0_count,
   input  [24:0] pre_instruction_source_in_stride0_max,
   input  [24:0] pre_instruction_source_in_stride0_min,
   input  [23:0] pre_instruction_source_in_stride1,
   input  [23:0] pre_instruction_source_in_stride1_count,
   input  [24:0] pre_instruction_source_in_stride1_max,
   input  [24:0] pre_instruction_source_in_stride1_min,
   input  [23:0] pre_instruction_source_in_stride2,
   input  [23:0] pre_instruction_source_in_stride2_count,
   input  [24:0] pre_instruction_source_in_stride2_max,
   input  [24:0] pre_instruction_source_in_stride2_min,
   input  [23:0] pre_instruction_source_in_stride3,
   input  [23:0] pre_instruction_source_in_stride3_count,
   input  [24:0] pre_instruction_source_in_stride3_max,
   input  [24:0] pre_instruction_source_in_stride3_min,
   input  [23:0] pre_instruction_source_in_stride4,
   input  [23:0] pre_instruction_source_in_stride4_count,
   input  [24:0] pre_instruction_source_in_stride4_max,
   input  [24:0] pre_instruction_source_in_stride4_min,
   input  [24:0] pre_instruction_source_in_burst_max,
   input  [24:0] pre_instruction_source_in_burst_max2,
   input  [24:0] pre_instruction_source_in_burst_max_init,
   input  [2:0] pre_instruction_source_in_burst_max_index,
   input  [24:0] pre_instruction_source_in_burst_min,
   input  [31:0] pre_instruction_source_in_bar,
   input  [23:0] pre_instruction_source_in_count,
   input  [23:0] pre_instruction_source_in_burststride,
   input  pre_instruction_source_in_double_precision,
   input  [1:0] pre_instruction_source_in_data_model,
   input  pre_instruction_source_in_scatter,
   input  [23:0] pre_instruction_source_in_totalcount,
   input  [5:0] pre_instruction_source_in_mcast,
   input  [15:0] pre_instruction_source_in_data,
   input  pre_instruction_source_in_repeat,
   input  [1:0] pre_instruction_source_in_datatype,
   input  [1:0] pre_instruction_source_in_bus_id,
   input  [23:0] pre_instruction_source_in_bufsize,
   input  [23:0] pre_instruction_source_in_burst_max_len,
   input  [23:0] pre_instruction_dest_in_stride0,
   input  [23:0] pre_instruction_dest_in_stride0_count,
   input  [24:0] pre_instruction_dest_in_stride0_max,
   input  [24:0] pre_instruction_dest_in_stride0_min,
   input  [23:0] pre_instruction_dest_in_stride1,
   input  [23:0] pre_instruction_dest_in_stride1_count,
   input  [24:0] pre_instruction_dest_in_stride1_max,
   input  [24:0] pre_instruction_dest_in_stride1_min,
   input  [23:0] pre_instruction_dest_in_stride2,
   input  [23:0] pre_instruction_dest_in_stride2_count,
   input  [24:0] pre_instruction_dest_in_stride2_max,
   input  [24:0] pre_instruction_dest_in_stride2_min,
   input  [23:0] pre_instruction_dest_in_stride3,
   input  [23:0] pre_instruction_dest_in_stride3_count,
   input  [24:0] pre_instruction_dest_in_stride3_max,
   input  [24:0] pre_instruction_dest_in_stride3_min,
   input  [23:0] pre_instruction_dest_in_stride4,
   input  [23:0] pre_instruction_dest_in_stride4_count,
   input  [24:0] pre_instruction_dest_in_stride4_max,
   input  [24:0] pre_instruction_dest_in_stride4_min,
   input  [24:0] pre_instruction_dest_in_burst_max,
   input  [24:0] pre_instruction_dest_in_burst_max2,
   input  [24:0] pre_instruction_dest_in_burst_max_init,
   input  [2:0] pre_instruction_dest_in_burst_max_index,
   input  [24:0] pre_instruction_dest_in_burst_min,
   input  [31:0] pre_instruction_dest_in_bar,
   input  [23:0] pre_instruction_dest_in_count,
   input  [23:0] pre_instruction_dest_in_burststride,
   input  pre_instruction_dest_in_double_precision,
   input  [1:0] pre_instruction_dest_in_data_model,
   input  pre_instruction_dest_in_scatter,
   input  [23:0] pre_instruction_dest_in_totalcount,
   input  [5:0] pre_instruction_dest_in_mcast,
   input  [15:0] pre_instruction_dest_in_data,
   input  pre_instruction_dest_in_repeat,
   input  [1:0] pre_instruction_dest_in_datatype,
   input  [1:0] pre_instruction_dest_in_bus_id,
   input  [23:0] pre_instruction_dest_in_bufsize,
   input  [23:0] pre_instruction_dest_in_burst_max_len,
   input  [1:0] pre_instruction_bus_id_source_in,
   input  [1:0] pre_instruction_bus_id_dest_in,
   input  instruction_source_addr_mode_in,
   input  instruction_dest_addr_mode_in,
   input  [1:0] instruction_bus_id_source_in,
   input  [1:0] instruction_data_type_source_in,
   input  [1:0] instruction_data_model_source_in,
   input  [1:0] instruction_bus_id_dest_in,
   input  [1:0] instruction_data_type_dest_in,
   input  [1:0] instruction_data_model_dest_in,
   input  [23:0] instruction_gen_len_in,
   input  [5:0] instruction_mcast_in,
   input  instruction_thread_in,
   input  [15:0] instruction_data_in,
   input  instruction_repeat_in,
   input  [14:0] wr_maxburstlen_in,
   input  [2:0] wr_full_in,
   input  [2:0] waitreq_in,
   input  [71:0] gen_bar_in,
   output ready_out,
   output [2:0] gen_valid_out,
   output gen_vm_out,
   output gen_fork_out,
   output [1:0] gen_data_flow_out,
   output gen_src_stream_out,
   output gen_dest_stream_out,
   output [1:0] gen_stream_id_out,
   output [2:0] gen_src_vector_out,
   output [2:0] gen_dst_vector_out,
   output [1:0] gen_src_scatter_out,
   output [1:0] gen_dst_scatter_out,
   output [3:0] gen_src_start_out,
   output [3:0] gen_src_end_out,
   output [3:0] gen_dst_end_out,
   output [31:0] gen_addr_source_out,
   output gen_addr_source_mode_out,
   output [31:0] gen_addr_dest_out,
   output gen_addr_dest_mode_out,
   output gen_eof_out,
   output [1:0] gen_bus_id_source_out,
   output [1:0] gen_data_type_source_out,
   output [1:0] gen_data_model_source_out,
   output [1:0] gen_bus_id_dest_out,
   output gen_busy_dest_out,
   output [1:0] gen_data_type_dest_out,
   output [1:0] gen_data_model_dest_out,
   output [4:0] gen_burstlen_source_out,
   output [4:0] gen_burstlen_dest_out,
   output gen_thread_out,
   output [5:0] gen_mcast_out,
   output [63:0] gen_data_out,
   output [31:0] log_out,
   output log_valid_out);
  wire [775:0] n26310_o;
  wire [775:0] n26311_o;
  wire [775:0] n26312_o;
  wire [775:0] n26313_o;
  wire [775:0] s_template_r;
  wire [23:0] s_i0_r;
  wire [23:0] s_i1_r;
  wire [23:0] s_i2_r;
  wire [23:0] s_i3_r;
  wire [23:0] s_i4_r;
  wire [23:0] s_i0_count_r;
  wire [23:0] s_i1_count_r;
  wire [23:0] s_i2_count_r;
  wire [23:0] s_i3_count_r;
  wire [23:0] s_i4_count_r;
  wire [23:0] s_burstlen_r;
  wire [23:0] s_burstpos_r;
  reg [23:0] s_burstremain_r;
  reg s_valid_r;
  wire [24:0] s_i0_start_r;
  wire [24:0] s_i1_start_r;
  wire [24:0] s_i2_start_r;
  wire [24:0] s_i3_start_r;
  wire [24:0] s_i4_start_r;
  wire [23:0] s_burstpos_stride_r;
  wire [24:0] s_burstpos_start_r;
  wire [3:0] s_burstpos_start_rr;
  wire [3:0] s_burstpos_start_rrr;
  wire [3:0] s_burstpos_start_rrrr;
  wire [26:0] s_burstpos_end_r;
  wire [3:0] s_burstpos_end_rr;
  wire [3:0] s_burstpos_end_rrr;
  wire [26:0] d_burstpos_end_r;
  wire [3:0] d_burstpos_end_rr;
  wire [3:0] d_burstpos_end_rrr;
  wire [775:0] d_template_r;
  wire [23:0] d_i0_r;
  wire [23:0] d_i1_r;
  wire [23:0] d_i2_r;
  wire [23:0] d_i3_r;
  wire [23:0] d_i4_r;
  wire [23:0] d_i0_count_r;
  wire [23:0] d_i1_count_r;
  wire [23:0] d_i2_count_r;
  wire [23:0] d_i3_count_r;
  wire [23:0] d_i4_count_r;
  wire [24:0] d_burst_max_r;
  wire [23:0] d_burstlen_r;
  wire [23:0] d_burstpos_r;
  reg [23:0] d_burstremain_r;
  reg d_valid_r;
  wire [23:0] currlen_r;
  wire [23:0] currlen_new;
  wire reload;
  wire s_burstlen_wrap;
  wire s_i0_wrap;
  wire s_i1_wrap;
  wire s_i2_wrap;
  wire s_i3_wrap;
  wire s_i4_wrap;
  wire [23:0] s_burstlen_new;
  wire [23:0] s_burstpos_new;
  wire [23:0] s_i0_new;
  wire [23:0] s_i1_new;
  wire [23:0] s_i2_new;
  wire [23:0] s_i3_new;
  wire [23:0] s_i4_new;
  wire [23:0] s_i0_count_new;
  wire [23:0] s_i1_count_new;
  wire [23:0] s_i2_count_new;
  wire [23:0] s_i3_count_new;
  wire [23:0] s_i4_count_new;
  wire [24:0] s_burstpos_start_new;
  wire [24:0] s_i0_start_new;
  wire [24:0] s_i1_start_new;
  wire [24:0] s_i2_start_new;
  wire [24:0] s_i3_start_new;
  wire [24:0] s_i4_start_new;
  wire d_burstlen_wrap;
  wire d_i0_wrap;
  wire d_i1_wrap;
  wire d_i2_wrap;
  wire d_i3_wrap;
  wire d_i4_wrap;
  wire [23:0] d_burstlen_new;
  wire [23:0] d_burstpos_new;
  wire [23:0] d_i0_new;
  wire [23:0] d_i1_new;
  wire [23:0] d_i2_new;
  wire [23:0] d_i3_new;
  wire [23:0] d_i4_new;
  wire [23:0] d_i0_new2;
  wire [23:0] d_i1_new2;
  wire [23:0] d_i2_new2;
  wire [23:0] d_i3_new2;
  wire [23:0] d_i4_new2;
  wire [23:0] d_i0_count_new;
  wire [23:0] d_i1_count_new;
  wire [23:0] d_i2_count_new;
  wire [23:0] d_i3_count_new;
  wire [23:0] d_i4_count_new;
  wire running_r;
  wire running_rr;
  wire running_rrr;
  wire running_rrrr;
  wire [2:0] gen_valid_r;
  wire [1:0] dp_dst_bus_id_r;
  wire [1:0] dp_dst_bus_id_rr;
  wire [1:0] dp_dst_bus_id_rrr;
  wire [1:0] dp_dst_bus_id_rrrr;
  wire [1:0] dp_src_bus_id_r;
  wire [1:0] dp_src_bus_id_rr;
  wire [1:0] dp_src_bus_id_rrr;
  wire [1:0] dp_src_bus_id_rrrr;
  wire [1:0] dp_dst_data_type_r;
  wire [1:0] dp_dst_data_type_rr;
  wire [1:0] dp_dst_data_type_rrr;
  wire [1:0] dp_dst_data_type_rrrr;
  wire [1:0] dp_src_data_type_r;
  wire [1:0] dp_src_data_type_rr;
  wire [1:0] dp_src_data_type_rrr;
  wire [1:0] dp_src_data_type_rrrr;
  wire [1:0] dp_src_data_model_r;
  wire [1:0] dp_src_data_model_rr;
  wire [1:0] dp_src_data_model_rrr;
  wire [1:0] dp_src_data_model_rrrr;
  wire [1:0] dp_dst_data_model_r;
  wire [1:0] dp_dst_data_model_rr;
  wire [1:0] dp_dst_data_model_rrr;
  wire [1:0] dp_dst_data_model_rrrr;
  wire dp_thread_r;
  wire dp_thread_rr;
  wire dp_thread_rrr;
  wire dp_thread_rrrr;
  reg [5:0] dp_mcast_r;
  reg [5:0] dp_mcast_rr;
  reg [5:0] dp_mcast_rrr;
  reg [5:0] dp_mcast_rrrr;
  wire [63:0] data_r;
  wire [63:0] data_rr;
  wire [63:0] data_rrr;
  wire [63:0] data_rrrr;
  wire [23:0] s_bufsize_r;
  wire [23:0] s_bufsize_rr;
  wire [23:0] s_temp1_r;
  wire [31:0] s_temp2_r;
  wire [23:0] s_temp3_r;
  wire [23:0] s_temp4_r;
  wire [23:0] s_temp5_r;
  wire [31:0] s_temp4_rr;
  wire [31:0] s_gen_addr_r;
  wire [4:0] s_gen_burstlen_r;
  wire [4:0] s_gen_burstlen_rr;
  wire s_gen_burstlen_progress_r;
  wire s_i0_valid;
  wire s_i1_valid;
  wire s_i2_valid;
  wire s_i3_valid;
  wire s_i4_valid;
  wire s_burst_valid;
  wire s_i0_start_valid;
  wire s_i1_start_valid;
  wire s_i2_start_valid;
  wire s_i3_start_valid;
  wire s_i4_start_valid;
  wire s_burst_start_valid;
  wire [23:0] d_bufsize_r;
  wire [23:0] d_bufsize_rr;
  wire [23:0] d_temp1_r;
  wire [31:0] d_temp2_r;
  wire [23:0] d_temp3_r;
  wire [23:0] d_temp4_r;
  wire [23:0] d_temp5_r;
  wire [31:0] d_temp4_rr;
  wire [31:0] d_gen_addr_r;
  wire [4:0] d_gen_burstlen_r;
  wire [4:0] d_gen_burstlen_rr;
  wire d_i0_valid;
  wire d_i1_valid;
  wire d_i2_valid;
  wire d_i3_valid;
  wire d_i4_valid;
  wire d_burst_valid;
  wire eof_r;
  wire eof_rr;
  wire eof_rrr;
  wire eof_rrrr;
  reg done_r;
  wire repeat_r;
  wire [1:0] data_flow_r;
  wire [1:0] data_flow_rr;
  wire [1:0] data_flow_rrr;
  wire [1:0] data_flow_rrrr;
  wire stream_src_r;
  wire stream_src_rr;
  wire stream_src_rrr;
  wire stream_src_rrrr;
  wire stream_dest_r;
  wire stream_dest_rr;
  wire stream_dest_rrr;
  wire stream_dest_rrrr;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire [1:0] stream_id_r;
  wire [1:0] stream_id_rr;
  wire [1:0] stream_id_rrr;
  wire [1:0] stream_id_rrrr;
  wire src_double_r;
  wire src_double_rr;
  wire src_double_rrr;
  wire dst_double_r;
  wire dst_double_rr;
  wire dst_double_rrr;
  wire [2:0] src_vector_r;
  wire [2:0] src_vector_rr;
  wire [2:0] src_vector_rrr;
  wire [2:0] src_vector_rrrr;
  wire [2:0] dst_vector_r;
  wire [2:0] dst_vector_rr;
  wire [2:0] dst_vector_rrr;
  wire [2:0] dst_vector_rrrr;
  wire src_addr_mode_r;
  wire src_addr_mode_rr;
  wire src_addr_mode_rrr;
  wire src_addr_mode_rrrr;
  wire dst_addr_mode_r;
  wire dst_addr_mode_rr;
  wire dst_addr_mode_rrr;
  wire dst_addr_mode_rrrr;
  wire [1:0] src_scatter_r;
  wire [1:0] src_scatter_rr;
  wire [1:0] src_scatter_rrr;
  wire [1:0] src_scatter_rrrr;
  wire [1:0] dst_scatter_r;
  wire [1:0] dst_scatter_rr;
  wire [1:0] dst_scatter_rrr;
  wire [1:0] dst_scatter_rrrr;
  wire [2:0] src_vector;
  wire [2:0] dst_vector;
  wire [1:0] src_scatter;
  wire [1:0] dst_scatter;
  wire src_is_burst_r;
  wire src_is_burst_rr;
  wire dst_is_burst_r;
  wire dst_is_burst_rr;
  wire [2:0] src_is_vector_r;
  wire [2:0] dst_is_vector_r;
  wire [5:0] src_is_scatter_r;
  wire [5:0] dst_is_scatter_r;
  wire [24:0] s_burst_actual_max_r;
  wire [31:0] log;
  wire [31:0] log_r;
  wire log_valid_r;
  wire source_double_precision;
  wire dest_double_precision;
  wire waitreq;
  wire ready;
  wire gen_busy_dest_r;
  wire n26356_o;
  wire n26358_o;
  wire n26359_o;
  wire n26361_o;
  wire n26363_o;
  wire n26364_o;
  wire n26367_o;
  wire n26368_o;
  wire n26369_o;
  wire n26370_o;
  wire n26371_o;
  wire n26372_o;
  wire n26373_o;
  wire n26374_o;
  wire n26375_o;
  wire n26378_o;
  wire n26379_o;
  wire n26380_o;
  wire [23:0] n26383_o;
  wire n26394_o;
  wire [2:0] n26396_o;
  wire n26398_o;
  wire n26400_o;
  wire n26401_o;
  wire n26402_o;
  wire n26403_o;
  wire [23:0] n26404_o;
  wire n26406_o;
  wire [23:0] n26408_o;
  wire n26410_o;
  wire [1:0] n26413_o;
  wire [1:0] n26414_o;
  wire [1:0] n26415_o;
  wire [2:0] n26416_o;
  wire n26418_o;
  wire n26420_o;
  wire n26421_o;
  wire n26422_o;
  wire n26423_o;
  wire [23:0] n26424_o;
  wire n26426_o;
  wire [23:0] n26427_o;
  wire n26429_o;
  wire [1:0] n26430_o;
  wire [1:0] n26431_o;
  wire [1:0] n26432_o;
  wire n26434_o;
  wire [23:0] n26435_o;
  wire n26437_o;
  wire [23:0] n26438_o;
  wire n26440_o;
  wire [2:0] n26441_o;
  wire n26443_o;
  wire n26444_o;
  wire n26445_o;
  wire n26448_o;
  wire [23:0] n26449_o;
  wire n26451_o;
  wire [2:0] n26452_o;
  wire n26454_o;
  wire [2:0] n26455_o;
  wire n26457_o;
  wire n26458_o;
  wire [2:0] n26459_o;
  wire n26461_o;
  wire n26462_o;
  wire [2:0] n26463_o;
  wire n26465_o;
  wire n26466_o;
  wire [2:0] n26467_o;
  wire n26469_o;
  wire n26470_o;
  wire [23:0] n26471_o;
  wire n26473_o;
  wire n26474_o;
  wire [2:0] n26475_o;
  wire n26477_o;
  wire n26478_o;
  wire [2:0] n26479_o;
  wire n26481_o;
  wire n26482_o;
  wire [2:0] n26483_o;
  wire n26485_o;
  wire n26486_o;
  wire n26487_o;
  wire n26490_o;
  wire n26491_o;
  wire n26493_o;
  wire [23:0] n26494_o;
  wire n26496_o;
  wire [23:0] n26497_o;
  wire n26499_o;
  wire [2:0] n26500_o;
  wire n26502_o;
  wire n26503_o;
  wire n26504_o;
  wire n26507_o;
  wire [23:0] n26508_o;
  wire n26510_o;
  wire [2:0] n26511_o;
  wire n26513_o;
  wire [2:0] n26514_o;
  wire n26516_o;
  wire n26517_o;
  wire [2:0] n26518_o;
  wire n26520_o;
  wire n26521_o;
  wire [2:0] n26522_o;
  wire n26524_o;
  wire n26525_o;
  wire [2:0] n26526_o;
  wire n26528_o;
  wire n26529_o;
  wire [23:0] n26530_o;
  wire n26532_o;
  wire n26533_o;
  wire [2:0] n26534_o;
  wire n26536_o;
  wire n26537_o;
  wire [2:0] n26538_o;
  wire n26540_o;
  wire n26541_o;
  wire [2:0] n26542_o;
  wire n26544_o;
  wire n26545_o;
  wire n26546_o;
  wire n26549_o;
  wire n26550_o;
  wire [1:0] n26551_o;
  wire n26553_o;
  wire n26555_o;
  wire n26556_o;
  wire n26557_o;
  wire n26558_o;
  wire [23:0] n26559_o;
  wire n26561_o;
  wire [23:0] n26562_o;
  wire n26564_o;
  wire [1:0] n26565_o;
  wire [1:0] n26566_o;
  wire [1:0] n26567_o;
  wire [1:0] n26568_o;
  wire n26570_o;
  wire n26572_o;
  wire n26573_o;
  wire n26574_o;
  wire n26575_o;
  wire [23:0] n26576_o;
  wire n26578_o;
  wire [23:0] n26579_o;
  wire n26581_o;
  wire [1:0] n26582_o;
  wire [1:0] n26583_o;
  wire [1:0] n26584_o;
  wire n26586_o;
  wire [23:0] n26587_o;
  wire n26589_o;
  wire [23:0] n26590_o;
  wire n26592_o;
  wire [1:0] n26593_o;
  wire n26595_o;
  wire n26596_o;
  wire n26597_o;
  wire n26600_o;
  wire [23:0] n26601_o;
  wire n26603_o;
  wire [1:0] n26604_o;
  wire n26606_o;
  wire [1:0] n26607_o;
  wire n26609_o;
  wire n26610_o;
  wire [1:0] n26611_o;
  wire n26613_o;
  wire n26614_o;
  wire [1:0] n26615_o;
  wire n26617_o;
  wire n26618_o;
  wire [1:0] n26619_o;
  wire n26621_o;
  wire n26622_o;
  wire [23:0] n26623_o;
  wire n26625_o;
  wire n26626_o;
  wire [1:0] n26627_o;
  wire n26629_o;
  wire n26630_o;
  wire [1:0] n26631_o;
  wire n26633_o;
  wire n26634_o;
  wire [1:0] n26635_o;
  wire n26637_o;
  wire n26638_o;
  wire n26639_o;
  wire n26642_o;
  wire n26643_o;
  wire n26645_o;
  wire [23:0] n26646_o;
  wire n26648_o;
  wire [23:0] n26649_o;
  wire n26651_o;
  wire [1:0] n26652_o;
  wire n26654_o;
  wire n26655_o;
  wire n26656_o;
  wire n26659_o;
  wire [23:0] n26660_o;
  wire n26662_o;
  wire [1:0] n26663_o;
  wire n26665_o;
  wire [1:0] n26666_o;
  wire n26668_o;
  wire n26669_o;
  wire [1:0] n26670_o;
  wire n26672_o;
  wire n26673_o;
  wire [1:0] n26674_o;
  wire n26676_o;
  wire n26677_o;
  wire [1:0] n26678_o;
  wire n26680_o;
  wire n26681_o;
  wire [23:0] n26682_o;
  wire n26684_o;
  wire n26685_o;
  wire [1:0] n26686_o;
  wire n26688_o;
  wire n26689_o;
  wire [1:0] n26690_o;
  wire n26692_o;
  wire n26693_o;
  wire [1:0] n26694_o;
  wire n26696_o;
  wire n26697_o;
  wire n26698_o;
  wire n26701_o;
  wire n26702_o;
  wire n26703_o;
  wire n26705_o;
  wire n26707_o;
  wire n26708_o;
  wire n26709_o;
  wire n26710_o;
  wire [23:0] n26711_o;
  wire n26713_o;
  wire [23:0] n26714_o;
  wire n26716_o;
  wire [1:0] n26717_o;
  wire [1:0] n26718_o;
  wire [1:0] n26719_o;
  wire n26720_o;
  wire n26722_o;
  wire n26724_o;
  wire n26725_o;
  wire n26726_o;
  wire n26727_o;
  wire [23:0] n26728_o;
  wire n26730_o;
  wire [23:0] n26731_o;
  wire n26733_o;
  wire [1:0] n26734_o;
  wire [1:0] n26735_o;
  wire [1:0] n26736_o;
  wire n26738_o;
  wire [23:0] n26739_o;
  wire n26741_o;
  wire [23:0] n26742_o;
  wire n26744_o;
  wire n26745_o;
  wire n26747_o;
  wire n26748_o;
  wire n26749_o;
  wire n26752_o;
  wire [23:0] n26753_o;
  wire n26755_o;
  wire n26756_o;
  wire n26758_o;
  wire n26759_o;
  wire n26761_o;
  wire n26762_o;
  wire n26763_o;
  wire n26765_o;
  wire n26766_o;
  wire n26767_o;
  wire n26769_o;
  wire n26770_o;
  wire n26771_o;
  wire n26773_o;
  wire n26774_o;
  wire [23:0] n26775_o;
  wire n26777_o;
  wire n26778_o;
  wire n26779_o;
  wire n26781_o;
  wire n26782_o;
  wire n26783_o;
  wire n26785_o;
  wire n26786_o;
  wire n26787_o;
  wire n26789_o;
  wire n26790_o;
  wire n26791_o;
  wire n26794_o;
  wire n26795_o;
  wire n26797_o;
  wire [23:0] n26798_o;
  wire n26800_o;
  wire [23:0] n26801_o;
  wire n26803_o;
  wire n26804_o;
  wire n26806_o;
  wire n26807_o;
  wire n26808_o;
  wire n26811_o;
  wire [23:0] n26812_o;
  wire n26814_o;
  wire n26815_o;
  wire n26817_o;
  wire n26818_o;
  wire n26820_o;
  wire n26821_o;
  wire n26822_o;
  wire n26824_o;
  wire n26825_o;
  wire n26826_o;
  wire n26828_o;
  wire n26829_o;
  wire n26830_o;
  wire n26832_o;
  wire n26833_o;
  wire [23:0] n26834_o;
  wire n26836_o;
  wire n26837_o;
  wire n26838_o;
  wire n26840_o;
  wire n26841_o;
  wire n26842_o;
  wire n26844_o;
  wire n26845_o;
  wire n26846_o;
  wire n26848_o;
  wire n26849_o;
  wire n26850_o;
  wire n26853_o;
  wire n26854_o;
  wire [2:0] n26855_o;
  wire [2:0] n26857_o;
  wire [5:0] n26859_o;
  wire [5:0] n26861_o;
  wire n26880_o;
  wire [1:0] n26881_o;
  wire n26883_o;
  wire n26884_o;
  wire n26885_o;
  wire n26886_o;
  wire n26887_o;
  wire n26888_o;
  wire [1:0] n26889_o;
  wire n26891_o;
  wire n26892_o;
  wire n26893_o;
  wire n26894_o;
  wire n26895_o;
  wire n26896_o;
  wire [1:0] n26897_o;
  wire [1:0] n26898_o;
  wire n26899_o;
  wire [1:0] n26900_o;
  wire n26902_o;
  wire n26903_o;
  wire n26904_o;
  wire [1:0] n26905_o;
  wire n26907_o;
  wire n26908_o;
  wire n26909_o;
  wire [1:0] n26910_o;
  wire [1:0] n26911_o;
  wire n26912_o;
  wire [1:0] n26913_o;
  wire n26915_o;
  wire n26916_o;
  wire n26917_o;
  wire [1:0] n26918_o;
  wire n26920_o;
  wire n26921_o;
  wire n26922_o;
  wire [1:0] n26923_o;
  wire [1:0] n26924_o;
  wire [2:0] n26927_o;
  wire [2:0] n26930_o;
  wire [1:0] n26932_o;
  wire [1:0] n26934_o;
  wire [2:0] n26936_o;
  wire [2:0] n26938_o;
  wire [1:0] n26939_o;
  wire [1:0] n26940_o;
  wire [2:0] n26942_o;
  wire [2:0] n26944_o;
  wire [1:0] n26945_o;
  wire [1:0] n26946_o;
  wire [23:0] n26949_o;
  wire [23:0] n26950_o;
  wire [23:0] n26951_o;
  wire [23:0] n26952_o;
  wire [23:0] n26953_o;
  wire [23:0] n26954_o;
  wire [23:0] n26955_o;
  wire [23:0] n26956_o;
  wire [23:0] n26957_o;
  wire [23:0] n26958_o;
  wire [23:0] n26959_o;
  wire [23:0] n26960_o;
  wire [23:0] n26961_o;
  wire [24:0] n26963_o;
  wire [24:0] n26964_o;
  wire [23:0] n26965_o;
  wire [24:0] n26967_o;
  wire [24:0] n26968_o;
  wire [23:0] n26969_o;
  wire [24:0] n26971_o;
  wire [24:0] n26972_o;
  wire [23:0] n26973_o;
  wire [24:0] n26975_o;
  wire [24:0] n26976_o;
  wire [23:0] n26977_o;
  wire [24:0] n26979_o;
  wire [24:0] n26980_o;
  wire [23:0] n26981_o;
  wire [24:0] n26983_o;
  wire [24:0] n26984_o;
  wire [23:0] n26986_o;
  wire [23:0] n26988_o;
  wire [23:0] n26990_o;
  wire [23:0] n26992_o;
  wire [23:0] n26994_o;
  wire [23:0] n26996_o;
  wire [23:0] n26997_o;
  wire [23:0] n26998_o;
  wire [23:0] n26999_o;
  wire [23:0] n27000_o;
  wire [23:0] n27001_o;
  wire [23:0] n27002_o;
  wire [23:0] n27003_o;
  wire [23:0] n27004_o;
  wire [23:0] n27005_o;
  wire [23:0] n27006_o;
  wire [23:0] n27007_o;
  wire [23:0] n27008_o;
  wire [22:0] n27009_o;
  wire [23:0] n27011_o;
  wire [23:0] n27012_o;
  wire [22:0] n27013_o;
  wire [23:0] n27015_o;
  wire [23:0] n27016_o;
  wire [22:0] n27017_o;
  wire [23:0] n27019_o;
  wire [23:0] n27020_o;
  wire [22:0] n27021_o;
  wire [23:0] n27023_o;
  wire [23:0] n27024_o;
  wire [22:0] n27025_o;
  wire [23:0] n27027_o;
  wire [23:0] n27028_o;
  wire [23:0] n27030_o;
  wire [23:0] n27032_o;
  wire [23:0] n27034_o;
  wire [23:0] n27036_o;
  wire [23:0] n27038_o;
  localparam n27039_o = 1'b0;
  wire n27041_o;
  wire n27042_o;
  wire n27043_o;
  wire [2:0] n27046_o;
  wire n27048_o;
  wire n27049_o;
  wire [23:0] n27052_o;
  wire n27053_o;
  wire n27054_o;
  wire [23:0] n27057_o;
  wire n27058_o;
  wire n27059_o;
  wire [23:0] n27062_o;
  wire n27063_o;
  wire n27064_o;
  wire [23:0] n27067_o;
  wire n27068_o;
  wire n27069_o;
  wire [23:0] n27072_o;
  wire n27073_o;
  wire n27074_o;
  wire [23:0] n27077_o;
  wire n27078_o;
  wire n27079_o;
  wire [23:0] n27082_o;
  wire n27083_o;
  wire n27084_o;
  wire n27085_o;
  wire n27086_o;
  wire n27087_o;
  wire [23:0] n27090_o;
  wire n27091_o;
  wire n27092_o;
  wire n27093_o;
  wire n27094_o;
  wire n27095_o;
  wire [23:0] n27098_o;
  wire n27099_o;
  wire n27100_o;
  wire n27101_o;
  wire n27102_o;
  wire n27103_o;
  wire [23:0] n27106_o;
  wire n27107_o;
  wire n27108_o;
  wire n27109_o;
  wire n27110_o;
  wire n27111_o;
  wire [23:0] n27114_o;
  wire n27115_o;
  wire n27116_o;
  wire n27117_o;
  wire n27118_o;
  wire n27119_o;
  wire [23:0] n27122_o;
  wire n27123_o;
  wire n27124_o;
  wire n27125_o;
  wire n27126_o;
  wire n27127_o;
  wire n27129_o;
  wire n27130_o;
  wire n27131_o;
  wire n27132_o;
  wire n27133_o;
  wire n27134_o;
  wire n27135_o;
  wire n27136_o;
  wire n27137_o;
  wire n27138_o;
  wire [24:0] n27140_o;
  wire [24:0] n27141_o;
  wire n27143_o;
  wire n27144_o;
  wire [23:0] n27147_o;
  wire n27148_o;
  wire n27149_o;
  wire [23:0] n27152_o;
  wire n27153_o;
  wire n27154_o;
  wire [23:0] n27157_o;
  wire n27158_o;
  wire n27159_o;
  wire [23:0] n27162_o;
  wire n27163_o;
  wire n27164_o;
  wire [23:0] n27167_o;
  wire n27168_o;
  wire n27169_o;
  wire [23:0] n27172_o;
  wire n27173_o;
  wire n27174_o;
  wire [23:0] n27177_o;
  wire n27178_o;
  wire n27179_o;
  wire n27180_o;
  wire n27181_o;
  wire n27182_o;
  wire [23:0] n27185_o;
  wire n27186_o;
  wire n27187_o;
  wire n27188_o;
  wire n27189_o;
  wire n27190_o;
  wire [23:0] n27193_o;
  wire n27194_o;
  wire n27195_o;
  wire n27196_o;
  wire n27197_o;
  wire n27198_o;
  wire [23:0] n27201_o;
  wire n27202_o;
  wire n27203_o;
  wire n27204_o;
  wire n27205_o;
  wire n27206_o;
  wire [23:0] n27209_o;
  wire n27210_o;
  wire n27211_o;
  wire n27212_o;
  wire n27213_o;
  wire n27214_o;
  wire [23:0] n27217_o;
  wire n27218_o;
  wire n27219_o;
  wire n27220_o;
  wire n27221_o;
  wire n27222_o;
  wire n27234_o;
  wire n27236_o;
  wire n27238_o;
  wire n27240_o;
  wire n27242_o;
  wire n27244_o;
  wire n27246_o;
  wire n27248_o;
  wire [23:0] n27252_o;
  wire [23:0] n27253_o;
  wire [23:0] n27254_o;
  wire [31:0] n27255_o;
  wire [23:0] n27256_o;
  wire [23:0] n27257_o;
  wire [23:0] n27258_o;
  wire [23:0] n27259_o;
  wire [23:0] n27260_o;
  wire [31:0] n27261_o;
  wire [31:0] n27262_o;
  wire [31:0] n27264_o;
  wire [31:0] n27265_o;
  wire n27269_o;
  wire [4:0] n27273_o;
  wire n27275_o;
  wire n27278_o;
  wire [26:0] n27279_o;
  wire [23:0] n27280_o;
  wire [26:0] n27281_o;
  wire [26:0] n27282_o;
  wire [26:0] n27284_o;
  wire [26:0] n27286_o;
  wire [26:0] n27287_o;
  wire n27288_o;
  wire [22:0] n27289_o;
  wire n27291_o;
  wire [3:0] n27292_o;
  wire [3:0] n27294_o;
  wire [3:0] n27296_o;
  wire [22:0] n27297_o;
  wire [24:0] n27298_o;
  wire [24:0] n27299_o;
  wire [24:0] n27300_o;
  wire [24:0] n27302_o;
  wire [24:0] n27303_o;
  wire n27305_o;
  wire [24:0] n27306_o;
  wire n27307_o;
  wire [3:0] n27308_o;
  wire [3:0] n27309_o;
  wire [3:0] n27311_o;
  wire [22:0] n27313_o;
  wire [23:0] n27315_o;
  wire [23:0] n27316_o;
  wire n27318_o;
  wire [22:0] n27319_o;
  wire n27322_o;
  wire [21:0] n27323_o;
  wire n27326_o;
  wire [20:0] n27327_o;
  wire [23:0] n27329_o;
  wire [23:0] n27330_o;
  wire [23:0] n27331_o;
  wire [23:0] n27332_o;
  wire [23:0] n27333_o;
  wire [23:0] n27334_o;
  wire n27335_o;
  wire n27336_o;
  wire n27337_o;
  wire n27338_o;
  wire n27339_o;
  wire n27340_o;
  wire n27341_o;
  wire n27342_o;
  wire n27343_o;
  wire n27344_o;
  wire n27345_o;
  wire n27346_o;
  wire n27348_o;
  wire [18:0] n27349_o;
  wire n27351_o;
  wire [4:0] n27352_o;
  wire n27354_o;
  wire n27355_o;
  wire [4:0] n27356_o;
  wire [4:0] n27358_o;
  wire n27359_o;
  wire [18:0] n27360_o;
  wire n27362_o;
  wire [4:0] n27363_o;
  wire n27364_o;
  wire n27365_o;
  wire [4:0] n27366_o;
  wire [4:0] n27368_o;
  wire [4:0] n27370_o;
  wire [4:0] n27371_o;
  wire [4:0] n27373_o;
  wire n27374_o;
  wire [4:0] n27377_o;
  wire [4:0] n27378_o;
  wire [4:0] n27381_o;
  wire [1:0] n27383_o;
  wire [2:0] n27385_o;
  wire [2:0] n27386_o;
  wire n27387_o;
  wire n27388_o;
  wire [21:0] n27389_o;
  wire n27391_o;
  wire [3:0] n27392_o;
  wire [3:0] n27395_o;
  wire [3:0] n27396_o;
  wire [3:0] n27398_o;
  wire [1:0] n27399_o;
  wire [2:0] n27401_o;
  wire [2:0] n27402_o;
  wire [23:0] n27403_o;
  wire [23:0] n27404_o;
  wire [23:0] n27405_o;
  wire [31:0] n27406_o;
  wire [23:0] n27407_o;
  wire [23:0] n27408_o;
  wire [23:0] n27409_o;
  wire [23:0] n27410_o;
  wire [23:0] n27411_o;
  wire [31:0] n27412_o;
  wire [31:0] n27413_o;
  wire [31:0] n27415_o;
  wire [31:0] n27416_o;
  wire [26:0] n27417_o;
  wire [23:0] n27418_o;
  wire [26:0] n27419_o;
  wire [26:0] n27420_o;
  wire [26:0] n27422_o;
  wire [26:0] n27424_o;
  wire [26:0] n27425_o;
  wire n27426_o;
  wire [22:0] n27427_o;
  wire n27429_o;
  wire [3:0] n27430_o;
  wire [3:0] n27432_o;
  wire [3:0] n27434_o;
  wire [22:0] n27435_o;
  wire [24:0] n27436_o;
  wire [24:0] n27437_o;
  wire [24:0] n27438_o;
  wire [24:0] n27440_o;
  wire [24:0] n27441_o;
  wire n27443_o;
  wire [24:0] n27444_o;
  wire n27445_o;
  wire [3:0] n27446_o;
  wire [3:0] n27447_o;
  wire [3:0] n27449_o;
  wire [22:0] n27451_o;
  wire [23:0] n27453_o;
  wire [23:0] n27454_o;
  wire n27456_o;
  wire [22:0] n27457_o;
  wire n27460_o;
  wire [21:0] n27461_o;
  wire n27464_o;
  wire [20:0] n27465_o;
  wire [23:0] n27467_o;
  wire [23:0] n27468_o;
  wire [23:0] n27469_o;
  wire [23:0] n27470_o;
  wire [23:0] n27471_o;
  wire [23:0] n27472_o;
  wire n27473_o;
  wire n27474_o;
  wire n27475_o;
  wire n27476_o;
  wire n27477_o;
  wire n27478_o;
  wire n27480_o;
  wire [18:0] n27481_o;
  wire n27483_o;
  wire [4:0] n27484_o;
  wire n27486_o;
  wire n27487_o;
  wire [4:0] n27488_o;
  wire [4:0] n27490_o;
  wire n27491_o;
  wire [18:0] n27492_o;
  wire n27494_o;
  wire [4:0] n27495_o;
  wire n27496_o;
  wire n27497_o;
  wire [4:0] n27498_o;
  wire [4:0] n27500_o;
  wire [4:0] n27502_o;
  wire [4:0] n27503_o;
  wire [4:0] n27505_o;
  wire n27506_o;
  wire [4:0] n27509_o;
  wire [4:0] n27510_o;
  wire [4:0] n27513_o;
  wire [2:0] n27536_o;
  wire n27632_o;
  reg [24:0] n28032_burst_min_v;
  wire n28038_o;
  wire n28040_o;
  wire n28041_o;
  wire n28042_o;
  wire n28046_o;
  wire [23:0] n28047_o;
  wire [23:0] n28048_o;
  wire [24:0] n28049_o;
  wire [24:0] n28050_o;
  wire [23:0] n28051_o;
  wire [23:0] n28052_o;
  wire [24:0] n28053_o;
  wire [24:0] n28054_o;
  wire [23:0] n28055_o;
  wire [23:0] n28056_o;
  wire [24:0] n28057_o;
  wire [24:0] n28058_o;
  wire [23:0] n28059_o;
  wire [23:0] n28060_o;
  wire [24:0] n28061_o;
  wire [24:0] n28062_o;
  wire [23:0] n28063_o;
  wire [23:0] n28064_o;
  wire [24:0] n28065_o;
  wire [24:0] n28066_o;
  wire [21:0] n28067_o;
  wire n28068_o;
  wire n28069_o;
  wire n28070_o;
  wire n28071_o;
  wire n28072_o;
  wire n28073_o;
  wire n28074_o;
  wire n28075_o;
  wire n28076_o;
  wire [24:0] n28077_o;
  wire [23:0] n28078_o;
  wire [31:0] n28079_o;
  wire [23:0] n28080_o;
  wire n28082_o;
  wire [20:0] n28083_o;
  wire n28086_o;
  wire [21:0] n28087_o;
  wire n28090_o;
  wire [22:0] n28091_o;
  wire [23:0] n28093_o;
  wire [23:0] n28094_o;
  wire [23:0] n28095_o;
  wire [23:0] n28096_o;
  wire [23:0] n28097_o;
  wire [23:0] n28098_o;
  wire [23:0] n28099_o;
  wire [24:0] n28100_o;
  wire [24:0] n28102_o;
  wire [24:0] n28103_o;
  wire [24:0] n28104_o;
  wire [23:0] n28105_o;
  wire n28107_o;
  wire n28110_o;
  wire n28112_o;
  wire [1:0] n28113_o;
  wire n28115_o;
  wire [1:0] n28116_o;
  wire n28118_o;
  wire [23:0] n28121_o;
  wire [23:0] n28123_o;
  wire n28125_o;
  wire [1:0] n28126_o;
  wire n28128_o;
  wire [1:0] n28129_o;
  wire n28131_o;
  wire [23:0] n28134_o;
  wire [23:0] n28136_o;
  wire n28138_o;
  wire [1:0] n28139_o;
  wire n28141_o;
  wire [1:0] n28142_o;
  wire n28144_o;
  wire [23:0] n28147_o;
  wire [23:0] n28149_o;
  wire [23:0] n28150_o;
  wire [23:0] n28151_o;
  wire [23:0] n28152_o;
  wire [23:0] n28153_o;
  wire [23:0] n28155_o;
  wire [23:0] n28156_o;
  wire [23:0] n28157_o;
  wire [23:0] n28158_o;
  wire [24:0] n28159_o;
  wire [23:0] n28160_o;
  wire [23:0] n28161_o;
  wire [24:0] n28162_o;
  wire [23:0] n28163_o;
  wire [23:0] n28164_o;
  wire [24:0] n28165_o;
  wire [23:0] n28166_o;
  wire [23:0] n28167_o;
  wire [24:0] n28168_o;
  wire [23:0] n28169_o;
  wire [23:0] n28170_o;
  wire [24:0] n28171_o;
  wire [31:0] n28172_o;
  wire [23:0] n28173_o;
  wire [24:0] n28174_o;
  wire [24:0] n28175_o;
  wire [24:0] n28176_o;
  wire [2:0] n28177_o;
  wire [23:0] n28178_o;
  wire n28180_o;
  wire [20:0] n28181_o;
  wire n28184_o;
  wire [21:0] n28185_o;
  wire n28188_o;
  wire [22:0] n28189_o;
  wire [23:0] n28191_o;
  wire [23:0] n28192_o;
  wire [23:0] n28193_o;
  wire [23:0] n28194_o;
  wire [23:0] n28195_o;
  wire [23:0] n28196_o;
  wire [23:0] n28197_o;
  wire [23:0] n28198_o;
  wire n28200_o;
  wire n28203_o;
  wire n28205_o;
  wire [1:0] n28206_o;
  wire n28208_o;
  wire [1:0] n28210_o;
  wire n28212_o;
  wire [23:0] n28215_o;
  wire [23:0] n28216_o;
  wire n28218_o;
  wire [1:0] n28219_o;
  wire n28221_o;
  wire [1:0] n28223_o;
  wire n28225_o;
  wire [23:0] n28228_o;
  wire [23:0] n28229_o;
  wire n28231_o;
  wire [1:0] n28232_o;
  wire n28234_o;
  wire [1:0] n28236_o;
  wire n28238_o;
  wire [23:0] n28241_o;
  wire [23:0] n28242_o;
  wire [23:0] n28243_o;
  wire [23:0] n28244_o;
  wire [23:0] n28245_o;
  wire [23:0] n28246_o;
  wire n28248_o;
  wire n28250_o;
  wire n28252_o;
  wire n28254_o;
  wire n28256_o;
  wire n28257_o;
  wire n28258_o;
  wire n28259_o;
  wire n28260_o;
  wire n28261_o;
  wire n28262_o;
  wire [1:0] n28265_o;
  wire n28266_o;
  wire n28267_o;
  wire n28268_o;
  wire n28269_o;
  wire [1:0] n28272_o;
  wire [1:0] n28274_o;
  wire [1:0] n28275_o;
  wire n28277_o;
  wire [20:0] n28279_o;
  wire [20:0] n28281_o;
  wire n28283_o;
  wire [21:0] n28285_o;
  wire [21:0] n28287_o;
  wire n28289_o;
  wire [22:0] n28291_o;
  wire [22:0] n28293_o;
  wire [23:0] n28295_o;
  wire [23:0] n28296_o;
  wire [23:0] n28297_o;
  wire [23:0] n28298_o;
  wire [23:0] n28299_o;
  wire [23:0] n28300_o;
  wire [23:0] n28301_o;
  wire n28303_o;
  wire n28306_o;
  wire [7:0] n28307_o;
  wire [7:0] n28308_o;
  wire [15:0] n28309_o;
  wire [7:0] n28310_o;
  wire [23:0] n28311_o;
  wire [7:0] n28312_o;
  wire [31:0] n28313_o;
  wire [7:0] n28314_o;
  wire [39:0] n28315_o;
  wire [7:0] n28316_o;
  wire [47:0] n28317_o;
  wire [7:0] n28318_o;
  wire [55:0] n28319_o;
  wire [7:0] n28320_o;
  wire [63:0] n28321_o;
  wire [7:0] n28322_o;
  wire [7:0] n28323_o;
  wire [15:0] n28324_o;
  wire [7:0] n28325_o;
  wire [23:0] n28326_o;
  wire [7:0] n28327_o;
  wire [31:0] n28328_o;
  wire [7:0] n28329_o;
  wire [39:0] n28330_o;
  wire [7:0] n28331_o;
  wire [47:0] n28332_o;
  wire [7:0] n28333_o;
  wire [55:0] n28334_o;
  wire [7:0] n28335_o;
  wire [63:0] n28336_o;
  wire [63:0] n28337_o;
  wire [23:0] n28338_o;
  wire n28340_o;
  wire n28343_o;
  wire [514:0] n28344_o;
  wire [104:0] n28345_o;
  wire [47:0] n28346_o;
  wire [72:0] n28354_o;
  wire [72:0] n28355_o;
  wire [72:0] n28356_o;
  wire [72:0] n28357_o;
  wire [72:0] n28358_o;
  wire [49:0] n28359_o;
  wire [79:0] n28360_o;
  wire [47:0] n28361_o;
  wire [24:0] n28380_o;
  wire [23:0] n28381_o;
  wire n28392_o;
  wire n28393_o;
  wire [24:0] n28411_o;
  wire [24:0] n28414_o;
  wire [24:0] n28415_o;
  wire [24:0] n28416_o;
  wire [24:0] n28417_o;
  wire [24:0] n28418_o;
  wire n28420_o;
  wire n28423_o;
  wire n28424_o;
  wire n28425_o;
  wire [24:0] n28426_o;
  wire n28427_o;
  wire [24:0] n28428_o;
  wire [24:0] n28429_o;
  wire n28430_o;
  wire [24:0] n28431_o;
  wire [24:0] n28432_o;
  wire [24:0] n28433_o;
  wire n28434_o;
  wire [24:0] n28435_o;
  wire [24:0] n28436_o;
  wire [24:0] n28437_o;
  wire [24:0] n28438_o;
  wire n28439_o;
  wire [24:0] n28440_o;
  wire [24:0] n28441_o;
  wire [24:0] n28442_o;
  wire [24:0] n28443_o;
  wire [24:0] n28444_o;
  wire n28445_o;
  wire [24:0] n28446_o;
  wire [24:0] n28447_o;
  wire [24:0] n28448_o;
  wire [24:0] n28449_o;
  wire [24:0] n28450_o;
  wire [24:0] n28451_o;
  wire [23:0] n28453_o;
  wire [23:0] n28455_o;
  wire [24:0] n28456_o;
  wire [24:0] n28457_o;
  wire [24:0] n28458_o;
  wire [24:0] n28459_o;
  wire [24:0] n28460_o;
  wire [24:0] n28461_o;
  wire n28462_o;
  wire [23:0] n28463_o;
  wire [23:0] n28465_o;
  wire [23:0] n28466_o;
  wire [23:0] n28468_o;
  wire [24:0] n28469_o;
  wire [24:0] n28470_o;
  wire [24:0] n28471_o;
  wire [24:0] n28472_o;
  wire [24:0] n28473_o;
  wire [24:0] n28474_o;
  wire n28475_o;
  wire [23:0] n28476_o;
  wire [23:0] n28477_o;
  wire [23:0] n28479_o;
  wire [23:0] n28480_o;
  wire [23:0] n28481_o;
  wire [23:0] n28483_o;
  wire [24:0] n28484_o;
  wire [24:0] n28485_o;
  wire [24:0] n28486_o;
  wire [24:0] n28487_o;
  wire [24:0] n28488_o;
  wire [24:0] n28489_o;
  wire n28490_o;
  wire [23:0] n28491_o;
  wire [23:0] n28492_o;
  wire [23:0] n28493_o;
  wire [23:0] n28495_o;
  wire [23:0] n28496_o;
  wire [23:0] n28497_o;
  wire [23:0] n28498_o;
  wire [23:0] n28500_o;
  wire [24:0] n28501_o;
  wire [24:0] n28502_o;
  wire [24:0] n28503_o;
  wire [24:0] n28504_o;
  wire [24:0] n28505_o;
  wire [24:0] n28506_o;
  wire n28507_o;
  wire [23:0] n28508_o;
  wire [23:0] n28509_o;
  wire [23:0] n28510_o;
  wire [23:0] n28511_o;
  wire [23:0] n28513_o;
  wire [23:0] n28514_o;
  wire [23:0] n28515_o;
  wire [23:0] n28516_o;
  wire [23:0] n28517_o;
  wire [23:0] n28519_o;
  wire [24:0] n28520_o;
  wire [24:0] n28521_o;
  wire [24:0] n28522_o;
  wire [24:0] n28523_o;
  wire [24:0] n28524_o;
  wire [24:0] n28525_o;
  wire n28526_o;
  wire [23:0] n28527_o;
  wire [23:0] n28528_o;
  wire [23:0] n28529_o;
  wire [23:0] n28530_o;
  wire [23:0] n28531_o;
  wire [23:0] n28532_o;
  wire [23:0] n28533_o;
  wire [23:0] n28534_o;
  wire [23:0] n28535_o;
  wire [23:0] n28536_o;
  wire [23:0] n28538_o;
  wire [23:0] n28540_o;
  wire [24:0] n28541_o;
  wire [24:0] n28542_o;
  wire [24:0] n28543_o;
  wire [24:0] n28544_o;
  wire [24:0] n28545_o;
  wire [24:0] n28546_o;
  wire n28547_o;
  wire n28548_o;
  wire n28549_o;
  wire [2:0] n28550_o;
  wire n28552_o;
  wire [23:0] n28553_o;
  wire n28554_o;
  wire n28555_o;
  wire [24:0] n28556_o;
  wire [24:0] n28557_o;
  wire [24:0] n28558_o;
  wire n28559_o;
  wire [2:0] n28561_o;
  wire n28563_o;
  wire [23:0] n28564_o;
  wire n28565_o;
  wire n28566_o;
  wire [24:0] n28567_o;
  wire [24:0] n28568_o;
  wire [24:0] n28569_o;
  wire n28570_o;
  wire [2:0] n28572_o;
  wire n28574_o;
  wire [23:0] n28575_o;
  wire n28576_o;
  wire n28577_o;
  wire [24:0] n28578_o;
  wire [24:0] n28579_o;
  wire [24:0] n28580_o;
  wire n28581_o;
  wire [2:0] n28583_o;
  wire n28585_o;
  wire [23:0] n28586_o;
  wire n28587_o;
  wire n28588_o;
  wire [24:0] n28589_o;
  wire [24:0] n28590_o;
  wire [24:0] n28591_o;
  wire n28592_o;
  wire [2:0] n28594_o;
  wire n28596_o;
  wire [23:0] n28597_o;
  wire n28598_o;
  wire n28599_o;
  wire [24:0] n28600_o;
  wire [24:0] n28601_o;
  wire [24:0] n28602_o;
  wire [23:0] n28605_o;
  wire [23:0] n28607_o;
  wire n28608_o;
  wire [23:0] n28609_o;
  wire [23:0] n28611_o;
  wire [23:0] n28612_o;
  wire [23:0] n28614_o;
  wire [24:0] n28615_o;
  wire [23:0] n28616_o;
  wire [23:0] n28617_o;
  wire [23:0] n28619_o;
  wire [23:0] n28620_o;
  wire [23:0] n28621_o;
  wire [23:0] n28623_o;
  wire [24:0] n28624_o;
  wire [23:0] n28625_o;
  wire [23:0] n28626_o;
  wire [23:0] n28627_o;
  wire [23:0] n28629_o;
  wire [23:0] n28630_o;
  wire [23:0] n28631_o;
  wire [23:0] n28632_o;
  wire [23:0] n28634_o;
  wire [24:0] n28635_o;
  wire [23:0] n28636_o;
  wire [23:0] n28637_o;
  wire [23:0] n28638_o;
  wire [23:0] n28639_o;
  wire [23:0] n28641_o;
  wire [23:0] n28642_o;
  wire [23:0] n28643_o;
  wire [23:0] n28644_o;
  wire [23:0] n28645_o;
  wire [23:0] n28647_o;
  wire [24:0] n28648_o;
  wire [23:0] n28649_o;
  wire [23:0] n28650_o;
  wire [23:0] n28651_o;
  wire [23:0] n28652_o;
  wire [23:0] n28653_o;
  wire [23:0] n28654_o;
  wire [23:0] n28655_o;
  wire [23:0] n28656_o;
  wire [23:0] n28657_o;
  wire [23:0] n28658_o;
  wire [24:0] n28659_o;
  wire [23:0] n28661_o;
  wire [23:0] n28663_o;
  wire n28665_o;
  wire n28667_o;
  wire n28669_o;
  wire [23:0] n28671_o;
  wire [23:0] n28673_o;
  wire [23:0] n28675_o;
  wire [23:0] n28677_o;
  wire [23:0] n28679_o;
  wire [23:0] n28681_o;
  wire [23:0] n28683_o;
  wire [23:0] n28685_o;
  wire [23:0] n28687_o;
  wire [23:0] n28689_o;
  wire [23:0] n28691_o;
  wire [23:0] n28693_o;
  wire [24:0] n28694_o;
  wire [24:0] n28695_o;
  wire [24:0] n28696_o;
  wire [24:0] n28697_o;
  wire [24:0] n28698_o;
  wire n28699_o;
  wire [24:0] n28700_o;
  wire n28702_o;
  wire n28704_o;
  wire n28706_o;
  wire n28708_o;
  wire n28710_o;
  wire n28712_o;
  wire n28714_o;
  wire n28716_o;
  wire n28718_o;
  wire [23:0] n28720_o;
  wire [23:0] n28722_o;
  wire [23:0] n28724_o;
  wire [23:0] n28726_o;
  wire [23:0] n28728_o;
  wire [23:0] n28730_o;
  wire [23:0] n28732_o;
  wire [23:0] n28734_o;
  wire [23:0] n28736_o;
  wire [23:0] n28738_o;
  wire [24:0] n28739_o;
  wire [23:0] n28741_o;
  wire [23:0] n28743_o;
  wire [23:0] n28744_o;
  wire n28747_o;
  wire n28748_o;
  wire n28749_o;
  wire n28750_o;
  wire n28751_o;
  wire n28752_o;
  wire n28753_o;
  wire n28754_o;
  wire n28755_o;
  wire n28756_o;
  wire n28757_o;
  wire n28758_o;
  wire n28759_o;
  wire n28760_o;
  wire n28761_o;
  wire n28762_o;
  wire n28763_o;
  wire n28764_o;
  wire n28765_o;
  wire n28766_o;
  wire n28767_o;
  wire n28768_o;
  wire n28769_o;
  wire n28770_o;
  wire n28771_o;
  wire n28772_o;
  wire n28773_o;
  wire n28774_o;
  wire n28775_o;
  wire n28777_o;
  wire n28782_o;
  wire n28784_o;
  wire n28786_o;
  wire n28804_o;
  wire n28807_o;
  wire n28809_o;
  wire n28811_o;
  wire n28813_o;
  wire n28815_o;
  wire n28817_o;
  wire n28819_o;
  wire n28821_o;
  wire n28823_o;
  wire n28839_o;
  wire n28840_o;
  wire n28841_o;
  wire n28842_o;
  wire n28843_o;
  wire n28844_o;
  wire n28845_o;
  wire n28846_o;
  wire n28847_o;
  wire n28848_o;
  wire n28851_o;
  wire n28852_o;
  wire n28853_o;
  wire n28854_o;
  wire n28855_o;
  wire n28856_o;
  wire n28857_o;
  wire n28858_o;
  wire n28859_o;
  wire n28860_o;
  wire n28861_o;
  wire n28862_o;
  wire n28863_o;
  wire n28864_o;
  wire n28865_o;
  wire n28866_o;
  wire n28867_o;
  wire n28868_o;
  wire n28870_o;
  wire n28872_o;
  wire n29125_o;
  wire n29126_o;
  wire [24:0] n29127_o;
  reg [24:0] n29128_q;
  wire n29137_o;
  wire n29138_o;
  wire [47:0] n29139_o;
  wire [47:0] n29140_o;
  reg [47:0] n29141_q;
  wire n29142_o;
  wire n29143_o;
  wire [104:0] n29144_o;
  wire [104:0] n29145_o;
  reg [104:0] n29146_q;
  wire n29147_o;
  wire n29148_o;
  wire [514:0] n29149_o;
  wire [514:0] n29150_o;
  reg [514:0] n29151_q;
  wire [775:0] n29154_o;
  wire [23:0] n29155_o;
  reg [23:0] n29156_q;
  wire [23:0] n29157_o;
  reg [23:0] n29158_q;
  wire [23:0] n29159_o;
  reg [23:0] n29160_q;
  wire [23:0] n29161_o;
  reg [23:0] n29162_q;
  wire [23:0] n29163_o;
  reg [23:0] n29164_q;
  wire [23:0] n29165_o;
  reg [23:0] n29166_q;
  wire [23:0] n29167_o;
  reg [23:0] n29168_q;
  wire [23:0] n29169_o;
  reg [23:0] n29170_q;
  wire [23:0] n29171_o;
  reg [23:0] n29172_q;
  wire [23:0] n29173_o;
  reg [23:0] n29174_q;
  wire [23:0] n29175_o;
  reg [23:0] n29176_q;
  wire [23:0] n29177_o;
  reg [23:0] n29178_q;
  wire [23:0] n29181_o;
  reg [23:0] n29182_q;
  wire n29183_o;
  reg n29184_q;
  wire [24:0] n29185_o;
  reg [24:0] n29186_q;
  wire [24:0] n29187_o;
  reg [24:0] n29188_q;
  wire [24:0] n29189_o;
  reg [24:0] n29190_q;
  wire [24:0] n29191_o;
  reg [24:0] n29192_q;
  wire [24:0] n29193_o;
  reg [24:0] n29194_q;
  wire [23:0] n29195_o;
  reg [23:0] n29196_q;
  wire [24:0] n29197_o;
  reg [24:0] n29198_q;
  wire [3:0] n29199_o;
  reg [3:0] n29200_q;
  wire [3:0] n29201_o;
  reg [3:0] n29202_q;
  wire [3:0] n29203_o;
  reg [3:0] n29204_q;
  wire [26:0] n29205_o;
  reg [26:0] n29206_q;
  wire [3:0] n29207_o;
  reg [3:0] n29208_q;
  wire [3:0] n29209_o;
  reg [3:0] n29210_q;
  wire [26:0] n29211_o;
  reg [26:0] n29212_q;
  wire [3:0] n29213_o;
  reg [3:0] n29214_q;
  wire [3:0] n29215_o;
  reg [3:0] n29216_q;
  wire n29217_o;
  wire n29218_o;
  wire [47:0] n29219_o;
  wire [47:0] n29220_o;
  reg [47:0] n29221_q;
  wire n29222_o;
  wire n29223_o;
  wire [79:0] n29224_o;
  wire [79:0] n29225_o;
  reg [79:0] n29226_q;
  wire n29227_o;
  wire n29228_o;
  wire [2:0] n29229_o;
  wire [2:0] n29230_o;
  reg [2:0] n29231_q;
  wire n29232_o;
  wire n29233_o;
  wire [49:0] n29234_o;
  wire [49:0] n29235_o;
  reg [49:0] n29236_q;
  wire n29237_o;
  wire n29238_o;
  wire [72:0] n29239_o;
  wire [72:0] n29240_o;
  reg [72:0] n29241_q;
  wire n29242_o;
  wire n29243_o;
  wire [72:0] n29244_o;
  wire [72:0] n29245_o;
  reg [72:0] n29246_q;
  wire n29247_o;
  wire n29248_o;
  wire [72:0] n29249_o;
  wire [72:0] n29250_o;
  reg [72:0] n29251_q;
  wire n29252_o;
  wire n29253_o;
  wire [72:0] n29254_o;
  wire [72:0] n29255_o;
  reg [72:0] n29256_q;
  wire n29257_o;
  wire n29258_o;
  wire [72:0] n29259_o;
  wire [72:0] n29260_o;
  reg [72:0] n29261_q;
  wire [775:0] n29270_o;
  wire [23:0] n29271_o;
  reg [23:0] n29272_q;
  wire [23:0] n29273_o;
  reg [23:0] n29274_q;
  wire [23:0] n29275_o;
  reg [23:0] n29276_q;
  wire [23:0] n29277_o;
  reg [23:0] n29278_q;
  wire [23:0] n29279_o;
  reg [23:0] n29280_q;
  wire [23:0] n29281_o;
  reg [23:0] n29282_q;
  wire [23:0] n29283_o;
  reg [23:0] n29284_q;
  wire [23:0] n29285_o;
  reg [23:0] n29286_q;
  wire [23:0] n29287_o;
  reg [23:0] n29288_q;
  wire [23:0] n29289_o;
  reg [23:0] n29290_q;
  wire [24:0] n29291_o;
  reg [24:0] n29292_q;
  wire [23:0] n29293_o;
  reg [23:0] n29294_q;
  wire [23:0] n29295_o;
  reg [23:0] n29296_q;
  wire [23:0] n29299_o;
  reg [23:0] n29300_q;
  wire n29301_o;
  reg n29302_q;
  wire [23:0] n29303_o;
  reg [23:0] n29304_q;
  wire n29307_o;
  reg n29308_q;
  wire n29309_o;
  reg n29310_q;
  wire n29311_o;
  reg n29312_q;
  wire n29313_o;
  reg n29314_q;
  wire [2:0] n29315_o;
  reg [2:0] n29316_q;
  wire [1:0] n29317_o;
  reg [1:0] n29318_q;
  wire [1:0] n29319_o;
  reg [1:0] n29320_q;
  wire [1:0] n29321_o;
  reg [1:0] n29322_q;
  wire [1:0] n29323_o;
  reg [1:0] n29324_q;
  wire [1:0] n29325_o;
  reg [1:0] n29326_q;
  wire [1:0] n29327_o;
  reg [1:0] n29328_q;
  wire [1:0] n29329_o;
  reg [1:0] n29330_q;
  wire [1:0] n29331_o;
  reg [1:0] n29332_q;
  wire [1:0] n29333_o;
  reg [1:0] n29334_q;
  wire [1:0] n29335_o;
  reg [1:0] n29336_q;
  wire [1:0] n29337_o;
  reg [1:0] n29338_q;
  wire [1:0] n29339_o;
  reg [1:0] n29340_q;
  wire [1:0] n29341_o;
  reg [1:0] n29342_q;
  wire [1:0] n29343_o;
  reg [1:0] n29344_q;
  wire [1:0] n29345_o;
  reg [1:0] n29346_q;
  wire [1:0] n29347_o;
  reg [1:0] n29348_q;
  wire [1:0] n29349_o;
  reg [1:0] n29350_q;
  wire [1:0] n29351_o;
  reg [1:0] n29352_q;
  wire [1:0] n29353_o;
  reg [1:0] n29354_q;
  wire [1:0] n29355_o;
  reg [1:0] n29356_q;
  wire [1:0] n29357_o;
  reg [1:0] n29358_q;
  wire [1:0] n29359_o;
  reg [1:0] n29360_q;
  wire [1:0] n29361_o;
  reg [1:0] n29362_q;
  wire [1:0] n29363_o;
  reg [1:0] n29364_q;
  wire n29365_o;
  reg n29366_q;
  wire n29367_o;
  reg n29368_q;
  wire n29369_o;
  reg n29370_q;
  wire n29371_o;
  reg n29372_q;
  wire [5:0] n29373_o;
  reg [5:0] n29374_q;
  wire [5:0] n29375_o;
  reg [5:0] n29376_q;
  wire [5:0] n29377_o;
  reg [5:0] n29378_q;
  wire [5:0] n29379_o;
  reg [5:0] n29380_q;
  wire [63:0] n29381_o;
  reg [63:0] n29382_q;
  wire [63:0] n29383_o;
  reg [63:0] n29384_q;
  wire [63:0] n29385_o;
  reg [63:0] n29386_q;
  wire [63:0] n29387_o;
  reg [63:0] n29388_q;
  wire [23:0] n29389_o;
  reg [23:0] n29390_q;
  wire [23:0] n29391_o;
  reg [23:0] n29392_q;
  wire [23:0] n29393_o;
  reg [23:0] n29394_q;
  wire [31:0] n29395_o;
  reg [31:0] n29396_q;
  wire [23:0] n29397_o;
  reg [23:0] n29398_q;
  wire [23:0] n29399_o;
  reg [23:0] n29400_q;
  wire [23:0] n29401_o;
  reg [23:0] n29402_q;
  wire [31:0] n29403_o;
  reg [31:0] n29404_q;
  wire [31:0] n29405_o;
  reg [31:0] n29406_q;
  wire [4:0] n29407_o;
  reg [4:0] n29408_q;
  wire [4:0] n29409_o;
  reg [4:0] n29410_q;
  wire n29411_o;
  reg n29412_q;
  wire [23:0] n29413_o;
  reg [23:0] n29414_q;
  wire [23:0] n29415_o;
  reg [23:0] n29416_q;
  wire [23:0] n29417_o;
  reg [23:0] n29418_q;
  wire [31:0] n29419_o;
  reg [31:0] n29420_q;
  wire [23:0] n29421_o;
  reg [23:0] n29422_q;
  wire [23:0] n29423_o;
  reg [23:0] n29424_q;
  wire [23:0] n29425_o;
  reg [23:0] n29426_q;
  wire [31:0] n29427_o;
  reg [31:0] n29428_q;
  wire [31:0] n29429_o;
  reg [31:0] n29430_q;
  wire [4:0] n29431_o;
  reg [4:0] n29432_q;
  wire [4:0] n29433_o;
  reg [4:0] n29434_q;
  wire n29435_o;
  reg n29436_q;
  wire n29437_o;
  reg n29438_q;
  wire n29439_o;
  reg n29440_q;
  wire n29441_o;
  reg n29442_q;
  wire n29443_o;
  reg n29444_q;
  wire n29445_o;
  reg n29446_q;
  wire [1:0] n29447_o;
  reg [1:0] n29448_q;
  wire [1:0] n29449_o;
  reg [1:0] n29450_q;
  wire [1:0] n29451_o;
  reg [1:0] n29452_q;
  wire [1:0] n29453_o;
  reg [1:0] n29454_q;
  wire n29455_o;
  reg n29456_q;
  wire n29457_o;
  reg n29458_q;
  wire n29459_o;
  reg n29460_q;
  wire n29461_o;
  reg n29462_q;
  wire n29463_o;
  reg n29464_q;
  wire n29465_o;
  reg n29466_q;
  wire n29467_o;
  reg n29468_q;
  wire n29469_o;
  reg n29470_q;
  wire n29471_o;
  reg n29472_q;
  wire n29473_o;
  reg n29474_q;
  wire n29475_o;
  reg n29476_q;
  wire n29477_o;
  reg n29478_q;
  wire [1:0] n29479_o;
  reg [1:0] n29480_q;
  wire [1:0] n29481_o;
  reg [1:0] n29482_q;
  wire [1:0] n29483_o;
  reg [1:0] n29484_q;
  wire [1:0] n29485_o;
  reg [1:0] n29486_q;
  wire n29487_o;
  reg n29488_q;
  wire n29489_o;
  reg n29490_q;
  wire n29491_o;
  reg n29492_q;
  wire n29495_o;
  reg n29496_q;
  wire n29497_o;
  reg n29498_q;
  wire n29499_o;
  reg n29500_q;
  wire [2:0] n29503_o;
  reg [2:0] n29504_q;
  wire [2:0] n29505_o;
  reg [2:0] n29506_q;
  wire [2:0] n29507_o;
  reg [2:0] n29508_q;
  wire [2:0] n29509_o;
  reg [2:0] n29510_q;
  wire [2:0] n29511_o;
  reg [2:0] n29512_q;
  wire [2:0] n29513_o;
  reg [2:0] n29514_q;
  wire [2:0] n29515_o;
  reg [2:0] n29516_q;
  wire [2:0] n29517_o;
  reg [2:0] n29518_q;
  wire n29519_o;
  reg n29520_q;
  wire n29521_o;
  reg n29522_q;
  wire n29523_o;
  reg n29524_q;
  wire n29525_o;
  reg n29526_q;
  wire n29527_o;
  reg n29528_q;
  wire n29529_o;
  reg n29530_q;
  wire n29531_o;
  reg n29532_q;
  wire n29533_o;
  reg n29534_q;
  wire [1:0] n29535_o;
  reg [1:0] n29536_q;
  wire [1:0] n29537_o;
  reg [1:0] n29538_q;
  wire [1:0] n29539_o;
  reg [1:0] n29540_q;
  wire [1:0] n29541_o;
  reg [1:0] n29542_q;
  wire [1:0] n29543_o;
  reg [1:0] n29544_q;
  wire [1:0] n29545_o;
  reg [1:0] n29546_q;
  wire [1:0] n29547_o;
  reg [1:0] n29548_q;
  wire [1:0] n29549_o;
  reg [1:0] n29550_q;
  wire n29551_o;
  reg n29552_q;
  wire n29553_o;
  reg n29554_q;
  wire n29555_o;
  reg n29556_q;
  wire n29557_o;
  reg n29558_q;
  reg [2:0] n29560_q;
  reg [2:0] n29561_q;
  reg [5:0] n29562_q;
  reg [5:0] n29563_q;
  wire [24:0] n29564_o;
  reg [24:0] n29565_q;
  wire [31:0] n29566_o;
  wire [31:0] n29567_o;
  reg [31:0] n29568_q;
  reg n29569_q;
  reg n29572_q;
  wire n29573_o;
  wire n29574_o;
  wire n29575_o;
  wire n29576_o;
  wire n29577_o;
  wire n29578_o;
  wire n29579_o;
  wire [4:0] n29580_o;
  wire [4:0] n29581_o;
  wire [4:0] n29582_o;
  wire n29583_o;
  wire [4:0] n29584_o;
  wire n29585_o;
  wire [4:0] n29586_o;
  wire [4:0] n29587_o;
  wire [4:0] n29588_o;
  wire [4:0] n29589_o;
  wire n29590_o;
  wire [4:0] n29591_o;
  wire n29592_o;
  wire [4:0] n29593_o;
  wire n29594_o;
  wire n29595_o;
  wire n29596_o;
  wire n29597_o;
  wire n29598_o;
  wire n29599_o;
  wire n29600_o;
  assign ready_out = ready;
  assign gen_valid_out = gen_valid_r;
  assign gen_vm_out = vm_rrrr;
  assign gen_fork_out = n27039_o;
  assign gen_data_flow_out = data_flow_rrrr;
  assign gen_src_stream_out = stream_src_rrrr;
  assign gen_dest_stream_out = stream_dest_rrrr;
  assign gen_stream_id_out = stream_id_rrrr;
  assign gen_src_vector_out = src_vector_rrrr;
  assign gen_dst_vector_out = dst_vector_rrrr;
  assign gen_src_scatter_out = src_scatter_rrrr;
  assign gen_dst_scatter_out = dst_scatter_rrrr;
  assign gen_src_start_out = s_burstpos_start_rrrr;
  assign gen_src_end_out = s_burstpos_end_rrr;
  assign gen_dst_end_out = d_burstpos_end_rrr;
  assign gen_addr_source_out = s_gen_addr_r;
  assign gen_addr_source_mode_out = src_addr_mode_rrrr;
  assign gen_addr_dest_out = d_gen_addr_r;
  assign gen_addr_dest_mode_out = dst_addr_mode_rrrr;
  assign gen_eof_out = n27043_o;
  assign gen_bus_id_source_out = dp_src_bus_id_rrrr;
  assign gen_data_type_source_out = dp_src_data_type_rrrr;
  assign gen_data_model_source_out = dp_src_data_model_rrrr;
  assign gen_bus_id_dest_out = dp_dst_bus_id_rrrr;
  assign gen_busy_dest_out = gen_busy_dest_r;
  assign gen_data_type_dest_out = dp_dst_data_type_rrrr;
  assign gen_data_model_dest_out = dp_dst_data_model_rrrr;
  assign gen_burstlen_source_out = s_gen_burstlen_rr;
  assign gen_burstlen_dest_out = d_gen_burstlen_rr;
  assign gen_thread_out = dp_thread_rrrr;
  assign gen_mcast_out = dp_mcast_rrrr;
  assign gen_data_out = data_rrrr;
  assign log_out = log_r;
  assign log_valid_out = log_valid_r;
  /* ../../HW/src/util/fifo.vhd:46:9  */
  assign n26310_o = {instruction_source_in_burst_max_len, instruction_source_in_bufsize, instruction_source_in_bus_id, instruction_source_in_datatype, instruction_source_in_repeat, instruction_source_in_data, instruction_source_in_mcast, instruction_source_in_totalcount, instruction_source_in_scatter, instruction_source_in_data_model, instruction_source_in_double_precision, instruction_source_in_burststride, instruction_source_in_count, instruction_source_in_bar, instruction_source_in_burst_min, instruction_source_in_burst_max_index, instruction_source_in_burst_max_init, instruction_source_in_burst_max2, instruction_source_in_burst_max, instruction_source_in_stride4_min, instruction_source_in_stride4_max, instruction_source_in_stride4_count, instruction_source_in_stride4, instruction_source_in_stride3_min, instruction_source_in_stride3_max, instruction_source_in_stride3_count, instruction_source_in_stride3, instruction_source_in_stride2_min, instruction_source_in_stride2_max, instruction_source_in_stride2_count, instruction_source_in_stride2, instruction_source_in_stride1_min, instruction_source_in_stride1_max, instruction_source_in_stride1_count, instruction_source_in_stride1, instruction_source_in_stride0_min, instruction_source_in_stride0_max, instruction_source_in_stride0_count, instruction_source_in_stride0};
  /* ../../HW/src/util/fifo.vhd:45:9  */
  assign n26311_o = {instruction_dest_in_burst_max_len, instruction_dest_in_bufsize, instruction_dest_in_bus_id, instruction_dest_in_datatype, instruction_dest_in_repeat, instruction_dest_in_data, instruction_dest_in_mcast, instruction_dest_in_totalcount, instruction_dest_in_scatter, instruction_dest_in_data_model, instruction_dest_in_double_precision, instruction_dest_in_burststride, instruction_dest_in_count, instruction_dest_in_bar, instruction_dest_in_burst_min, instruction_dest_in_burst_max_index, instruction_dest_in_burst_max_init, instruction_dest_in_burst_max2, instruction_dest_in_burst_max, instruction_dest_in_stride4_min, instruction_dest_in_stride4_max, instruction_dest_in_stride4_count, instruction_dest_in_stride4, instruction_dest_in_stride3_min, instruction_dest_in_stride3_max, instruction_dest_in_stride3_count, instruction_dest_in_stride3, instruction_dest_in_stride2_min, instruction_dest_in_stride2_max, instruction_dest_in_stride2_count, instruction_dest_in_stride2, instruction_dest_in_stride1_min, instruction_dest_in_stride1_max, instruction_dest_in_stride1_count, instruction_dest_in_stride1, instruction_dest_in_stride0_min, instruction_dest_in_stride0_max, instruction_dest_in_stride0_count, instruction_dest_in_stride0};
  /* ../../HW/src/util/fifo.vhd:44:9  */
  assign n26312_o = {pre_instruction_source_in_burst_max_len, pre_instruction_source_in_bufsize, pre_instruction_source_in_bus_id, pre_instruction_source_in_datatype, pre_instruction_source_in_repeat, pre_instruction_source_in_data, pre_instruction_source_in_mcast, pre_instruction_source_in_totalcount, pre_instruction_source_in_scatter, pre_instruction_source_in_data_model, pre_instruction_source_in_double_precision, pre_instruction_source_in_burststride, pre_instruction_source_in_count, pre_instruction_source_in_bar, pre_instruction_source_in_burst_min, pre_instruction_source_in_burst_max_index, pre_instruction_source_in_burst_max_init, pre_instruction_source_in_burst_max2, pre_instruction_source_in_burst_max, pre_instruction_source_in_stride4_min, pre_instruction_source_in_stride4_max, pre_instruction_source_in_stride4_count, pre_instruction_source_in_stride4, pre_instruction_source_in_stride3_min, pre_instruction_source_in_stride3_max, pre_instruction_source_in_stride3_count, pre_instruction_source_in_stride3, pre_instruction_source_in_stride2_min, pre_instruction_source_in_stride2_max, pre_instruction_source_in_stride2_count, pre_instruction_source_in_stride2, pre_instruction_source_in_stride1_min, pre_instruction_source_in_stride1_max, pre_instruction_source_in_stride1_count, pre_instruction_source_in_stride1, pre_instruction_source_in_stride0_min, pre_instruction_source_in_stride0_max, pre_instruction_source_in_stride0_count, pre_instruction_source_in_stride0};
  /* ../../HW/src/util/fifo.vhd:43:9  */
  assign n26313_o = {pre_instruction_dest_in_burst_max_len, pre_instruction_dest_in_bufsize, pre_instruction_dest_in_bus_id, pre_instruction_dest_in_datatype, pre_instruction_dest_in_repeat, pre_instruction_dest_in_data, pre_instruction_dest_in_mcast, pre_instruction_dest_in_totalcount, pre_instruction_dest_in_scatter, pre_instruction_dest_in_data_model, pre_instruction_dest_in_double_precision, pre_instruction_dest_in_burststride, pre_instruction_dest_in_count, pre_instruction_dest_in_bar, pre_instruction_dest_in_burst_min, pre_instruction_dest_in_burst_max_index, pre_instruction_dest_in_burst_max_init, pre_instruction_dest_in_burst_max2, pre_instruction_dest_in_burst_max, pre_instruction_dest_in_stride4_min, pre_instruction_dest_in_stride4_max, pre_instruction_dest_in_stride4_count, pre_instruction_dest_in_stride4, pre_instruction_dest_in_stride3_min, pre_instruction_dest_in_stride3_max, pre_instruction_dest_in_stride3_count, pre_instruction_dest_in_stride3, pre_instruction_dest_in_stride2_min, pre_instruction_dest_in_stride2_max, pre_instruction_dest_in_stride2_count, pre_instruction_dest_in_stride2, pre_instruction_dest_in_stride1_min, pre_instruction_dest_in_stride1_max, pre_instruction_dest_in_stride1_count, pre_instruction_dest_in_stride1, pre_instruction_dest_in_stride0_min, pre_instruction_dest_in_stride0_max, pre_instruction_dest_in_stride0_count, pre_instruction_dest_in_stride0};
  /* ../../HW/src/dp/dp_gen.vhd:130:8  */
  assign s_template_r = n29154_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:131:8  */
  assign s_i0_r = n29156_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:132:8  */
  assign s_i1_r = n29158_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:133:8  */
  assign s_i2_r = n29160_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:134:8  */
  assign s_i3_r = n29162_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:135:8  */
  assign s_i4_r = n29164_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:136:8  */
  assign s_i0_count_r = n29166_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:137:8  */
  assign s_i1_count_r = n29168_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:138:8  */
  assign s_i2_count_r = n29170_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:139:8  */
  assign s_i3_count_r = n29172_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:140:8  */
  assign s_i4_count_r = n29174_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:141:8  */
  assign s_burstlen_r = n29176_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:142:8  */
  assign s_burstpos_r = n29178_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:144:8  */
  always @*
    s_burstremain_r = n29182_q; // (isignal)
  initial
    s_burstremain_r = 24'b111111111111111111111111;
  /* ../../HW/src/dp/dp_gen.vhd:145:8  */
  always @*
    s_valid_r = n29184_q; // (isignal)
  initial
    s_valid_r = 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:147:8  */
  assign s_i0_start_r = n29186_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:148:8  */
  assign s_i1_start_r = n29188_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:149:8  */
  assign s_i2_start_r = n29190_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:150:8  */
  assign s_i3_start_r = n29192_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:151:8  */
  assign s_i4_start_r = n29194_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:153:8  */
  assign s_burstpos_stride_r = n29196_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:154:8  */
  assign s_burstpos_start_r = n29198_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:155:8  */
  assign s_burstpos_start_rr = n29200_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:156:8  */
  assign s_burstpos_start_rrr = n29202_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:157:8  */
  assign s_burstpos_start_rrrr = n29204_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:159:8  */
  assign s_burstpos_end_r = n29206_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:160:8  */
  assign s_burstpos_end_rr = n29208_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:161:8  */
  assign s_burstpos_end_rrr = n29210_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:163:8  */
  assign d_burstpos_end_r = n29212_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:164:8  */
  assign d_burstpos_end_rr = n29214_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:165:8  */
  assign d_burstpos_end_rrr = n29216_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:168:8  */
  assign d_template_r = n29270_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:169:8  */
  assign d_i0_r = n29272_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:170:8  */
  assign d_i1_r = n29274_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:171:8  */
  assign d_i2_r = n29276_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:172:8  */
  assign d_i3_r = n29278_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:173:8  */
  assign d_i4_r = n29280_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:174:8  */
  assign d_i0_count_r = n29282_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:175:8  */
  assign d_i1_count_r = n29284_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:176:8  */
  assign d_i2_count_r = n29286_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:177:8  */
  assign d_i3_count_r = n29288_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:178:8  */
  assign d_i4_count_r = n29290_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:179:8  */
  assign d_burst_max_r = n29292_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:180:8  */
  assign d_burstlen_r = n29294_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:181:8  */
  assign d_burstpos_r = n29296_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:183:8  */
  always @*
    d_burstremain_r = n29300_q; // (isignal)
  initial
    d_burstremain_r = 24'b111111111111111111111111;
  /* ../../HW/src/dp/dp_gen.vhd:184:8  */
  always @*
    d_valid_r = n29302_q; // (isignal)
  initial
    d_valid_r = 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:186:8  */
  assign currlen_r = n29304_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:187:8  */
  assign currlen_new = n26383_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:189:8  */
  assign reload = n26380_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:191:8  */
  assign s_burstlen_wrap = n27054_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:192:8  */
  assign s_i0_wrap = n27059_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:193:8  */
  assign s_i1_wrap = n27064_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:194:8  */
  assign s_i2_wrap = n27069_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:195:8  */
  assign s_i3_wrap = n27074_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:196:8  */
  assign s_i4_wrap = n27079_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:197:8  */
  assign s_burstlen_new = n26949_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:198:8  */
  assign s_burstpos_new = n26951_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:199:8  */
  assign s_i0_new = n26953_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:200:8  */
  assign s_i1_new = n26955_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:201:8  */
  assign s_i2_new = n26957_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:202:8  */
  assign s_i3_new = n26959_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:203:8  */
  assign s_i4_new = n26961_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:204:8  */
  assign s_i0_count_new = n26986_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:205:8  */
  assign s_i1_count_new = n26988_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:206:8  */
  assign s_i2_count_new = n26990_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:207:8  */
  assign s_i3_count_new = n26992_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:208:8  */
  assign s_i4_count_new = n26994_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:210:8  */
  assign s_burstpos_start_new = n26964_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:211:8  */
  assign s_i0_start_new = n26968_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:212:8  */
  assign s_i1_start_new = n26972_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:213:8  */
  assign s_i2_start_new = n26976_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:214:8  */
  assign s_i3_start_new = n26980_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:215:8  */
  assign s_i4_start_new = n26984_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:217:8  */
  assign d_burstlen_wrap = n27149_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:218:8  */
  assign d_i0_wrap = n27154_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:219:8  */
  assign d_i1_wrap = n27159_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:220:8  */
  assign d_i2_wrap = n27164_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:221:8  */
  assign d_i3_wrap = n27169_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:222:8  */
  assign d_i4_wrap = n27174_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:223:8  */
  assign d_burstlen_new = n26996_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:224:8  */
  assign d_burstpos_new = n26998_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:225:8  */
  assign d_i0_new = n27000_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:226:8  */
  assign d_i1_new = n27002_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:227:8  */
  assign d_i2_new = n27004_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:228:8  */
  assign d_i3_new = n27006_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:229:8  */
  assign d_i4_new = n27008_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:230:8  */
  assign d_i0_new2 = n27012_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:231:8  */
  assign d_i1_new2 = n27016_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:232:8  */
  assign d_i2_new2 = n27020_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:233:8  */
  assign d_i3_new2 = n27024_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:234:8  */
  assign d_i4_new2 = n27028_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:235:8  */
  assign d_i0_count_new = n27030_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:236:8  */
  assign d_i1_count_new = n27032_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:237:8  */
  assign d_i2_count_new = n27034_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:238:8  */
  assign d_i3_count_new = n27036_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:239:8  */
  assign d_i4_count_new = n27038_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:241:8  */
  assign running_r = n29308_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:242:8  */
  assign running_rr = n29310_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:243:8  */
  assign running_rrr = n29312_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:244:8  */
  assign running_rrrr = n29314_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:245:8  */
  assign gen_valid_r = n29316_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:246:8  */
  assign dp_dst_bus_id_r = n29318_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:247:8  */
  assign dp_dst_bus_id_rr = n29320_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:248:8  */
  assign dp_dst_bus_id_rrr = n29322_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:249:8  */
  assign dp_dst_bus_id_rrrr = n29324_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:250:8  */
  assign dp_src_bus_id_r = n29326_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:251:8  */
  assign dp_src_bus_id_rr = n29328_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:252:8  */
  assign dp_src_bus_id_rrr = n29330_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:253:8  */
  assign dp_src_bus_id_rrrr = n29332_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:254:8  */
  assign dp_dst_data_type_r = n29334_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:255:8  */
  assign dp_dst_data_type_rr = n29336_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:256:8  */
  assign dp_dst_data_type_rrr = n29338_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:257:8  */
  assign dp_dst_data_type_rrrr = n29340_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:258:8  */
  assign dp_src_data_type_r = n29342_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:259:8  */
  assign dp_src_data_type_rr = n29344_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:260:8  */
  assign dp_src_data_type_rrr = n29346_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:261:8  */
  assign dp_src_data_type_rrrr = n29348_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:262:8  */
  assign dp_src_data_model_r = n29350_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:263:8  */
  assign dp_src_data_model_rr = n29352_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:264:8  */
  assign dp_src_data_model_rrr = n29354_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:265:8  */
  assign dp_src_data_model_rrrr = n29356_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:266:8  */
  assign dp_dst_data_model_r = n29358_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:267:8  */
  assign dp_dst_data_model_rr = n29360_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:268:8  */
  assign dp_dst_data_model_rrr = n29362_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:269:8  */
  assign dp_dst_data_model_rrrr = n29364_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:270:8  */
  assign dp_thread_r = n29366_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:271:8  */
  assign dp_thread_rr = n29368_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:272:8  */
  assign dp_thread_rrr = n29370_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:273:8  */
  assign dp_thread_rrrr = n29372_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:274:8  */
  always @*
    dp_mcast_r = n29374_q; // (isignal)
  initial
    dp_mcast_r = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:275:8  */
  always @*
    dp_mcast_rr = n29376_q; // (isignal)
  initial
    dp_mcast_rr = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:276:8  */
  always @*
    dp_mcast_rrr = n29378_q; // (isignal)
  initial
    dp_mcast_rrr = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:277:8  */
  always @*
    dp_mcast_rrrr = n29380_q; // (isignal)
  initial
    dp_mcast_rrrr = 6'b111111;
  /* ../../HW/src/dp/dp_gen.vhd:278:8  */
  assign data_r = n29382_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:279:8  */
  assign data_rr = n29384_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:280:8  */
  assign data_rrr = n29386_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:281:8  */
  assign data_rrrr = n29388_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:283:8  */
  assign s_bufsize_r = n29390_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:284:8  */
  assign s_bufsize_rr = n29392_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:285:8  */
  assign s_temp1_r = n29394_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:286:8  */
  assign s_temp2_r = n29396_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:287:8  */
  assign s_temp3_r = n29398_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:288:8  */
  assign s_temp4_r = n29400_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:289:8  */
  assign s_temp5_r = n29402_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:290:8  */
  assign s_temp4_rr = n29404_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:291:8  */
  assign s_gen_addr_r = n29406_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:292:8  */
  assign s_gen_burstlen_r = n29408_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:293:8  */
  assign s_gen_burstlen_rr = n29410_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:294:8  */
  assign s_gen_burstlen_progress_r = n29412_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:296:8  */
  assign s_i0_valid = n27087_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:297:8  */
  assign s_i1_valid = n27095_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:298:8  */
  assign s_i2_valid = n27103_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:299:8  */
  assign s_i3_valid = n27111_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:300:8  */
  assign s_i4_valid = n27119_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:301:8  */
  assign s_burst_valid = n27127_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:303:8  */
  assign s_i0_start_valid = n27130_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:304:8  */
  assign s_i1_start_valid = n27132_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:305:8  */
  assign s_i2_start_valid = n27134_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:306:8  */
  assign s_i3_start_valid = n27136_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:307:8  */
  assign s_i4_start_valid = n27138_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:308:8  */
  assign s_burst_start_valid = n27144_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:310:8  */
  assign d_bufsize_r = n29414_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:311:8  */
  assign d_bufsize_rr = n29416_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:312:8  */
  assign d_temp1_r = n29418_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:313:8  */
  assign d_temp2_r = n29420_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:314:8  */
  assign d_temp3_r = n29422_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:315:8  */
  assign d_temp4_r = n29424_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:316:8  */
  assign d_temp5_r = n29426_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:317:8  */
  assign d_temp4_rr = n29428_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:318:8  */
  assign d_gen_addr_r = n29430_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:319:8  */
  assign d_gen_burstlen_r = n29432_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:320:8  */
  assign d_gen_burstlen_rr = n29434_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:322:8  */
  assign d_i0_valid = n27182_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:323:8  */
  assign d_i1_valid = n27190_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:324:8  */
  assign d_i2_valid = n27198_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:325:8  */
  assign d_i3_valid = n27206_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:326:8  */
  assign d_i4_valid = n27214_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:327:8  */
  assign d_burst_valid = n27222_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:329:8  */
  assign eof_r = n29436_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:330:8  */
  assign eof_rr = n29438_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:331:8  */
  assign eof_rrr = n29440_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:332:8  */
  assign eof_rrrr = n29442_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:333:8  */
  always @*
    done_r = n29444_q; // (isignal)
  initial
    done_r = 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:335:8  */
  assign repeat_r = n29446_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:337:8  */
  assign data_flow_r = n29448_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:338:8  */
  assign data_flow_rr = n29450_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:339:8  */
  assign data_flow_rrr = n29452_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:340:8  */
  assign data_flow_rrrr = n29454_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:342:8  */
  assign stream_src_r = n29456_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:343:8  */
  assign stream_src_rr = n29458_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:344:8  */
  assign stream_src_rrr = n29460_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:345:8  */
  assign stream_src_rrrr = n29462_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:347:8  */
  assign stream_dest_r = n29464_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:348:8  */
  assign stream_dest_rr = n29466_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:349:8  */
  assign stream_dest_rrr = n29468_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:350:8  */
  assign stream_dest_rrrr = n29470_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:352:8  */
  assign vm_r = n29472_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:353:8  */
  assign vm_rr = n29474_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:354:8  */
  assign vm_rrr = n29476_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:355:8  */
  assign vm_rrrr = n29478_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:357:8  */
  assign stream_id_r = n29480_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:358:8  */
  assign stream_id_rr = n29482_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:359:8  */
  assign stream_id_rrr = n29484_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:360:8  */
  assign stream_id_rrrr = n29486_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:362:8  */
  assign src_double_r = n29488_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:363:8  */
  assign src_double_rr = n29490_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:364:8  */
  assign src_double_rrr = n29492_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:367:8  */
  assign dst_double_r = n29496_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:368:8  */
  assign dst_double_rr = n29498_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:369:8  */
  assign dst_double_rrr = n29500_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:372:8  */
  assign src_vector_r = n29504_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:373:8  */
  assign src_vector_rr = n29506_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:374:8  */
  assign src_vector_rrr = n29508_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:375:8  */
  assign src_vector_rrrr = n29510_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:377:8  */
  assign dst_vector_r = n29512_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:378:8  */
  assign dst_vector_rr = n29514_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:379:8  */
  assign dst_vector_rrr = n29516_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:380:8  */
  assign dst_vector_rrrr = n29518_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:382:8  */
  assign src_addr_mode_r = n29520_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:383:8  */
  assign src_addr_mode_rr = n29522_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:384:8  */
  assign src_addr_mode_rrr = n29524_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:385:8  */
  assign src_addr_mode_rrrr = n29526_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:387:8  */
  assign dst_addr_mode_r = n29528_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:388:8  */
  assign dst_addr_mode_rr = n29530_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:389:8  */
  assign dst_addr_mode_rrr = n29532_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:390:8  */
  assign dst_addr_mode_rrrr = n29534_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:392:8  */
  assign src_scatter_r = n29536_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:393:8  */
  assign src_scatter_rr = n29538_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:394:8  */
  assign src_scatter_rrr = n29540_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:395:8  */
  assign src_scatter_rrrr = n29542_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:397:8  */
  assign dst_scatter_r = n29544_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:398:8  */
  assign dst_scatter_rr = n29546_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:399:8  */
  assign dst_scatter_rrr = n29548_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:400:8  */
  assign dst_scatter_rrrr = n29550_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:402:8  */
  assign src_vector = n26942_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:403:8  */
  assign dst_vector = n26944_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:404:8  */
  assign src_scatter = n26945_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:405:8  */
  assign dst_scatter = n26946_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:407:8  */
  assign src_is_burst_r = n29552_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:408:8  */
  assign src_is_burst_rr = n29554_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:409:8  */
  assign dst_is_burst_r = n29556_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:410:8  */
  assign dst_is_burst_rr = n29558_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:413:8  */
  assign src_is_vector_r = n29560_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:414:8  */
  assign dst_is_vector_r = n29561_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:415:8  */
  assign src_is_scatter_r = n29562_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:416:8  */
  assign dst_is_scatter_r = n29563_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:418:8  */
  assign s_burst_actual_max_r = n29565_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:420:8  */
  assign log = n29566_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:421:8  */
  assign log_r = n29568_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:422:8  */
  assign log_valid_r = n29569_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:424:8  */
  assign source_double_precision = n26359_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:425:8  */
  assign dest_double_precision = n26364_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:427:8  */
  assign waitreq = n27049_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:429:8  */
  assign ready = n26375_o; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:441:8  */
  assign gen_busy_dest_r = n29572_q; // (signal)
  /* ../../HW/src/dp/dp_gen.vhd:452:50  */
  assign n26356_o = n26310_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:452:100  */
  assign n26358_o = instruction_bus_id_source_in != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:452:67  */
  assign n26359_o = n26358_o ? n26356_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:453:46  */
  assign n26361_o = n26311_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:453:94  */
  assign n26363_o = instruction_bus_id_dest_in != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:453:63  */
  assign n26364_o = n26363_o ? n26361_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:456:29  */
  assign n26367_o = ~running_r;
  /* ../../HW/src/dp/dp_gen.vhd:456:48  */
  assign n26368_o = ~running_rr;
  /* ../../HW/src/dp/dp_gen.vhd:456:34  */
  assign n26369_o = n26368_o & n26367_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:68  */
  assign n26370_o = ~running_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:456:53  */
  assign n26371_o = n26370_o & n26369_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:89  */
  assign n26372_o = ~running_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:456:73  */
  assign n26373_o = n26372_o & n26371_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:95  */
  assign n26374_o = reload & n26373_o;
  /* ../../HW/src/dp/dp_gen.vhd:456:14  */
  assign n26375_o = n26374_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:459:30  */
  assign n26378_o = ~running_r;
  /* ../../HW/src/dp/dp_gen.vhd:459:35  */
  assign n26379_o = n26378_o | done_r;
  /* ../../HW/src/dp/dp_gen.vhd:459:15  */
  assign n26380_o = n26379_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:462:25  */
  assign n26383_o = currlen_r - 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:531:12  */
  assign n26394_o = ~reset_in;
  /* ../../HW/src/dp/dp_gen.vhd:541:42  */
  assign n26396_o = n26312_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:541:62  */
  assign n26398_o = n26396_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:542:43  */
  assign n26400_o = pre_instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:541:98  */
  assign n26401_o = n26400_o & n26398_o;
  /* ../../HW/src/dp/dp_gen.vhd:543:37  */
  assign n26402_o = n26312_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:542:98  */
  assign n26403_o = n26402_o & n26401_o;
  /* ../../HW/src/dp/dp_gen.vhd:544:39  */
  assign n26404_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:544:50  */
  assign n26406_o = n26404_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:546:42  */
  assign n26408_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:546:53  */
  assign n26410_o = n26408_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:546:10  */
  assign n26413_o = n26410_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:544:10  */
  assign n26414_o = n26406_o ? 2'b01 : n26413_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:7  */
  assign n26415_o = n26403_o ? n26414_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:40  */
  assign n26416_o = n26313_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:555:60  */
  assign n26418_o = n26416_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:556:41  */
  assign n26420_o = pre_instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:96  */
  assign n26421_o = n26420_o & n26418_o;
  /* ../../HW/src/dp/dp_gen.vhd:557:35  */
  assign n26422_o = n26313_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:556:96  */
  assign n26423_o = n26422_o & n26421_o;
  /* ../../HW/src/dp/dp_gen.vhd:558:37  */
  assign n26424_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:558:48  */
  assign n26426_o = n26424_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:560:40  */
  assign n26427_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:560:51  */
  assign n26429_o = n26427_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:560:10  */
  assign n26430_o = n26429_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:558:10  */
  assign n26431_o = n26426_o ? 2'b01 : n26430_o;
  /* ../../HW/src/dp/dp_gen.vhd:555:7  */
  assign n26432_o = n26423_o ? n26431_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:569:42  */
  assign n26434_o = pre_instruction_bus_id_source_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:570:39  */
  assign n26435_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:570:50  */
  assign n26437_o = n26435_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:571:39  */
  assign n26438_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:571:50  */
  assign n26440_o = n26438_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:572:44  */
  assign n26441_o = n26312_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:572:64  */
  assign n26443_o = n26441_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:571:111  */
  assign n26444_o = n26443_o & n26440_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:111  */
  assign n26445_o = n26437_o | n26444_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:10  */
  assign n26448_o = n26445_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:577:39  */
  assign n26449_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:577:50  */
  assign n26451_o = n26449_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:578:46  */
  assign n26452_o = n26312_o[2:0];
  /* ../../HW/src/dp/dp_gen.vhd:578:66  */
  assign n26454_o = n26452_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:579:46  */
  assign n26455_o = n26312_o[100:98];
  /* ../../HW/src/dp/dp_gen.vhd:579:66  */
  assign n26457_o = n26455_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:578:90  */
  assign n26458_o = n26457_o & n26454_o;
  /* ../../HW/src/dp/dp_gen.vhd:580:46  */
  assign n26459_o = n26312_o[198:196];
  /* ../../HW/src/dp/dp_gen.vhd:580:66  */
  assign n26461_o = n26459_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:579:90  */
  assign n26462_o = n26461_o & n26458_o;
  /* ../../HW/src/dp/dp_gen.vhd:581:46  */
  assign n26463_o = n26312_o[296:294];
  /* ../../HW/src/dp/dp_gen.vhd:581:66  */
  assign n26465_o = n26463_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:580:90  */
  assign n26466_o = n26465_o & n26462_o;
  /* ../../HW/src/dp/dp_gen.vhd:582:46  */
  assign n26467_o = n26312_o[394:392];
  /* ../../HW/src/dp/dp_gen.vhd:582:66  */
  assign n26469_o = n26467_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:581:90  */
  assign n26470_o = n26469_o & n26466_o;
  /* ../../HW/src/dp/dp_gen.vhd:583:39  */
  assign n26471_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:583:50  */
  assign n26473_o = n26471_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:582:90  */
  assign n26474_o = n26473_o & n26470_o;
  /* ../../HW/src/dp/dp_gen.vhd:584:44  */
  assign n26475_o = n26312_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:584:64  */
  assign n26477_o = n26475_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:583:111  */
  assign n26478_o = n26477_o & n26474_o;
  /* ../../HW/src/dp/dp_gen.vhd:585:48  */
  assign n26479_o = n26312_o[492:490];
  /* ../../HW/src/dp/dp_gen.vhd:585:68  */
  assign n26481_o = n26479_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:584:99  */
  assign n26482_o = n26481_o & n26478_o;
  /* ../../HW/src/dp/dp_gen.vhd:586:42  */
  assign n26483_o = n26312_o[595:593];
  /* ../../HW/src/dp/dp_gen.vhd:586:62  */
  assign n26485_o = n26483_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:585:103  */
  assign n26486_o = n26485_o & n26482_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:111  */
  assign n26487_o = n26451_o | n26486_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:7  */
  assign n26490_o = n26487_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:569:7  */
  assign n26491_o = n26434_o ? n26448_o : n26490_o;
  /* ../../HW/src/dp/dp_gen.vhd:593:41  */
  assign n26493_o = pre_instruction_bus_id_dest_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:594:38  */
  assign n26494_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:594:49  */
  assign n26496_o = n26494_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:595:38  */
  assign n26497_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:595:49  */
  assign n26499_o = n26497_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:596:43  */
  assign n26500_o = n26313_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:596:63  */
  assign n26502_o = n26500_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:595:108  */
  assign n26503_o = n26502_o & n26499_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:108  */
  assign n26504_o = n26496_o | n26503_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:11  */
  assign n26507_o = n26504_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:601:35  */
  assign n26508_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:601:46  */
  assign n26510_o = n26508_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:602:42  */
  assign n26511_o = n26313_o[2:0];
  /* ../../HW/src/dp/dp_gen.vhd:602:62  */
  assign n26513_o = n26511_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:603:42  */
  assign n26514_o = n26313_o[100:98];
  /* ../../HW/src/dp/dp_gen.vhd:603:62  */
  assign n26516_o = n26514_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:602:86  */
  assign n26517_o = n26516_o & n26513_o;
  /* ../../HW/src/dp/dp_gen.vhd:604:42  */
  assign n26518_o = n26313_o[198:196];
  /* ../../HW/src/dp/dp_gen.vhd:604:62  */
  assign n26520_o = n26518_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:603:86  */
  assign n26521_o = n26520_o & n26517_o;
  /* ../../HW/src/dp/dp_gen.vhd:605:42  */
  assign n26522_o = n26313_o[296:294];
  /* ../../HW/src/dp/dp_gen.vhd:605:62  */
  assign n26524_o = n26522_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:604:86  */
  assign n26525_o = n26524_o & n26521_o;
  /* ../../HW/src/dp/dp_gen.vhd:606:42  */
  assign n26526_o = n26313_o[394:392];
  /* ../../HW/src/dp/dp_gen.vhd:606:62  */
  assign n26528_o = n26526_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:605:86  */
  assign n26529_o = n26528_o & n26525_o;
  /* ../../HW/src/dp/dp_gen.vhd:607:35  */
  assign n26530_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:607:46  */
  assign n26532_o = n26530_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:606:86  */
  assign n26533_o = n26532_o & n26529_o;
  /* ../../HW/src/dp/dp_gen.vhd:608:40  */
  assign n26534_o = n26313_o[627:625];
  /* ../../HW/src/dp/dp_gen.vhd:608:60  */
  assign n26536_o = n26534_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:607:105  */
  assign n26537_o = n26536_o & n26533_o;
  /* ../../HW/src/dp/dp_gen.vhd:609:44  */
  assign n26538_o = n26313_o[492:490];
  /* ../../HW/src/dp/dp_gen.vhd:609:64  */
  assign n26540_o = n26538_o == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:608:95  */
  assign n26541_o = n26540_o & n26537_o;
  /* ../../HW/src/dp/dp_gen.vhd:610:38  */
  assign n26542_o = n26313_o[595:593];
  /* ../../HW/src/dp/dp_gen.vhd:610:58  */
  assign n26544_o = n26542_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:609:99  */
  assign n26545_o = n26544_o & n26541_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:105  */
  assign n26546_o = n26510_o | n26545_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:5  */
  assign n26549_o = n26546_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:593:8  */
  assign n26550_o = n26493_o ? n26507_o : n26549_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:42  */
  assign n26551_o = n26312_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:541:62  */
  assign n26553_o = n26551_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:542:43  */
  assign n26555_o = pre_instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:541:98  */
  assign n26556_o = n26555_o & n26553_o;
  /* ../../HW/src/dp/dp_gen.vhd:543:37  */
  assign n26557_o = n26312_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:542:98  */
  assign n26558_o = n26557_o & n26556_o;
  /* ../../HW/src/dp/dp_gen.vhd:544:39  */
  assign n26559_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:544:50  */
  assign n26561_o = n26559_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:546:42  */
  assign n26562_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:546:53  */
  assign n26564_o = n26562_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:546:10  */
  assign n26565_o = n26564_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:544:10  */
  assign n26566_o = n26561_o ? 2'b01 : n26565_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:7  */
  assign n26567_o = n26558_o ? n26566_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:40  */
  assign n26568_o = n26313_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:555:60  */
  assign n26570_o = n26568_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:556:41  */
  assign n26572_o = pre_instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:96  */
  assign n26573_o = n26572_o & n26570_o;
  /* ../../HW/src/dp/dp_gen.vhd:557:35  */
  assign n26574_o = n26313_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:556:96  */
  assign n26575_o = n26574_o & n26573_o;
  /* ../../HW/src/dp/dp_gen.vhd:558:37  */
  assign n26576_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:558:48  */
  assign n26578_o = n26576_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:560:40  */
  assign n26579_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:560:51  */
  assign n26581_o = n26579_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:560:10  */
  assign n26582_o = n26581_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:558:10  */
  assign n26583_o = n26578_o ? 2'b01 : n26582_o;
  /* ../../HW/src/dp/dp_gen.vhd:555:7  */
  assign n26584_o = n26575_o ? n26583_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:569:42  */
  assign n26586_o = pre_instruction_bus_id_source_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:570:39  */
  assign n26587_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:570:50  */
  assign n26589_o = n26587_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:571:39  */
  assign n26590_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:571:50  */
  assign n26592_o = n26590_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:572:44  */
  assign n26593_o = n26312_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:572:64  */
  assign n26595_o = n26593_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:571:111  */
  assign n26596_o = n26595_o & n26592_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:111  */
  assign n26597_o = n26589_o | n26596_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:10  */
  assign n26600_o = n26597_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:577:39  */
  assign n26601_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:577:50  */
  assign n26603_o = n26601_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:578:46  */
  assign n26604_o = n26312_o[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:578:66  */
  assign n26606_o = n26604_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:579:46  */
  assign n26607_o = n26312_o[99:98];
  /* ../../HW/src/dp/dp_gen.vhd:579:66  */
  assign n26609_o = n26607_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:578:90  */
  assign n26610_o = n26609_o & n26606_o;
  /* ../../HW/src/dp/dp_gen.vhd:580:46  */
  assign n26611_o = n26312_o[197:196];
  /* ../../HW/src/dp/dp_gen.vhd:580:66  */
  assign n26613_o = n26611_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:579:90  */
  assign n26614_o = n26613_o & n26610_o;
  /* ../../HW/src/dp/dp_gen.vhd:581:46  */
  assign n26615_o = n26312_o[295:294];
  /* ../../HW/src/dp/dp_gen.vhd:581:66  */
  assign n26617_o = n26615_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:580:90  */
  assign n26618_o = n26617_o & n26614_o;
  /* ../../HW/src/dp/dp_gen.vhd:582:46  */
  assign n26619_o = n26312_o[393:392];
  /* ../../HW/src/dp/dp_gen.vhd:582:66  */
  assign n26621_o = n26619_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:581:90  */
  assign n26622_o = n26621_o & n26618_o;
  /* ../../HW/src/dp/dp_gen.vhd:583:39  */
  assign n26623_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:583:50  */
  assign n26625_o = n26623_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:582:90  */
  assign n26626_o = n26625_o & n26622_o;
  /* ../../HW/src/dp/dp_gen.vhd:584:44  */
  assign n26627_o = n26312_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:584:64  */
  assign n26629_o = n26627_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:583:111  */
  assign n26630_o = n26629_o & n26626_o;
  /* ../../HW/src/dp/dp_gen.vhd:585:48  */
  assign n26631_o = n26312_o[491:490];
  /* ../../HW/src/dp/dp_gen.vhd:585:68  */
  assign n26633_o = n26631_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:584:99  */
  assign n26634_o = n26633_o & n26630_o;
  /* ../../HW/src/dp/dp_gen.vhd:586:42  */
  assign n26635_o = n26312_o[594:593];
  /* ../../HW/src/dp/dp_gen.vhd:586:62  */
  assign n26637_o = n26635_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:585:103  */
  assign n26638_o = n26637_o & n26634_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:111  */
  assign n26639_o = n26603_o | n26638_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:7  */
  assign n26642_o = n26639_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:569:7  */
  assign n26643_o = n26586_o ? n26600_o : n26642_o;
  /* ../../HW/src/dp/dp_gen.vhd:593:41  */
  assign n26645_o = pre_instruction_bus_id_dest_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:594:38  */
  assign n26646_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:594:49  */
  assign n26648_o = n26646_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:595:38  */
  assign n26649_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:595:49  */
  assign n26651_o = n26649_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:596:43  */
  assign n26652_o = n26313_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:596:63  */
  assign n26654_o = n26652_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:595:108  */
  assign n26655_o = n26654_o & n26651_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:108  */
  assign n26656_o = n26648_o | n26655_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:11  */
  assign n26659_o = n26656_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:601:35  */
  assign n26660_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:601:46  */
  assign n26662_o = n26660_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:602:42  */
  assign n26663_o = n26313_o[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:602:62  */
  assign n26665_o = n26663_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:603:42  */
  assign n26666_o = n26313_o[99:98];
  /* ../../HW/src/dp/dp_gen.vhd:603:62  */
  assign n26668_o = n26666_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:602:86  */
  assign n26669_o = n26668_o & n26665_o;
  /* ../../HW/src/dp/dp_gen.vhd:604:42  */
  assign n26670_o = n26313_o[197:196];
  /* ../../HW/src/dp/dp_gen.vhd:604:62  */
  assign n26672_o = n26670_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:603:86  */
  assign n26673_o = n26672_o & n26669_o;
  /* ../../HW/src/dp/dp_gen.vhd:605:42  */
  assign n26674_o = n26313_o[295:294];
  /* ../../HW/src/dp/dp_gen.vhd:605:62  */
  assign n26676_o = n26674_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:604:86  */
  assign n26677_o = n26676_o & n26673_o;
  /* ../../HW/src/dp/dp_gen.vhd:606:42  */
  assign n26678_o = n26313_o[393:392];
  /* ../../HW/src/dp/dp_gen.vhd:606:62  */
  assign n26680_o = n26678_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:605:86  */
  assign n26681_o = n26680_o & n26677_o;
  /* ../../HW/src/dp/dp_gen.vhd:607:35  */
  assign n26682_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:607:46  */
  assign n26684_o = n26682_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:606:86  */
  assign n26685_o = n26684_o & n26681_o;
  /* ../../HW/src/dp/dp_gen.vhd:608:40  */
  assign n26686_o = n26313_o[626:625];
  /* ../../HW/src/dp/dp_gen.vhd:608:60  */
  assign n26688_o = n26686_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:607:105  */
  assign n26689_o = n26688_o & n26685_o;
  /* ../../HW/src/dp/dp_gen.vhd:609:44  */
  assign n26690_o = n26313_o[491:490];
  /* ../../HW/src/dp/dp_gen.vhd:609:64  */
  assign n26692_o = n26690_o == 2'b11;
  /* ../../HW/src/dp/dp_gen.vhd:608:95  */
  assign n26693_o = n26692_o & n26689_o;
  /* ../../HW/src/dp/dp_gen.vhd:610:38  */
  assign n26694_o = n26313_o[594:593];
  /* ../../HW/src/dp/dp_gen.vhd:610:58  */
  assign n26696_o = n26694_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:609:99  */
  assign n26697_o = n26696_o & n26693_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:105  */
  assign n26698_o = n26662_o | n26697_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:5  */
  assign n26701_o = n26698_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:593:8  */
  assign n26702_o = n26645_o ? n26659_o : n26701_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:42  */
  assign n26703_o = n26312_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:541:62  */
  assign n26705_o = n26703_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:542:43  */
  assign n26707_o = pre_instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:541:98  */
  assign n26708_o = n26707_o & n26705_o;
  /* ../../HW/src/dp/dp_gen.vhd:543:37  */
  assign n26709_o = n26312_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:542:98  */
  assign n26710_o = n26709_o & n26708_o;
  /* ../../HW/src/dp/dp_gen.vhd:544:39  */
  assign n26711_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:544:50  */
  assign n26713_o = n26711_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:546:42  */
  assign n26714_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:546:53  */
  assign n26716_o = n26714_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:546:10  */
  assign n26717_o = n26716_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:544:10  */
  assign n26718_o = n26713_o ? 2'b01 : n26717_o;
  /* ../../HW/src/dp/dp_gen.vhd:541:7  */
  assign n26719_o = n26710_o ? n26718_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:40  */
  assign n26720_o = n26313_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:555:60  */
  assign n26722_o = n26720_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:556:41  */
  assign n26724_o = pre_instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:555:96  */
  assign n26725_o = n26724_o & n26722_o;
  /* ../../HW/src/dp/dp_gen.vhd:557:35  */
  assign n26726_o = n26313_o[676];
  /* ../../HW/src/dp/dp_gen.vhd:556:96  */
  assign n26727_o = n26726_o & n26725_o;
  /* ../../HW/src/dp/dp_gen.vhd:558:37  */
  assign n26728_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:558:48  */
  assign n26730_o = n26728_o == 24'b000000000000000000001000;
  /* ../../HW/src/dp/dp_gen.vhd:560:40  */
  assign n26731_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:560:51  */
  assign n26733_o = n26731_o == 24'b000000000000000100000000;
  /* ../../HW/src/dp/dp_gen.vhd:560:10  */
  assign n26734_o = n26733_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:558:10  */
  assign n26735_o = n26730_o ? 2'b01 : n26734_o;
  /* ../../HW/src/dp/dp_gen.vhd:555:7  */
  assign n26736_o = n26727_o ? n26735_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:569:42  */
  assign n26738_o = pre_instruction_bus_id_source_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:570:39  */
  assign n26739_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:570:50  */
  assign n26741_o = n26739_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:571:39  */
  assign n26742_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:571:50  */
  assign n26744_o = n26742_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:572:44  */
  assign n26745_o = n26312_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:572:64  */
  assign n26747_o = n26745_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:571:111  */
  assign n26748_o = n26747_o & n26744_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:111  */
  assign n26749_o = n26741_o | n26748_o;
  /* ../../HW/src/dp/dp_gen.vhd:570:10  */
  assign n26752_o = n26749_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:577:39  */
  assign n26753_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:577:50  */
  assign n26755_o = n26753_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:578:46  */
  assign n26756_o = n26312_o[0];
  /* ../../HW/src/dp/dp_gen.vhd:578:66  */
  assign n26758_o = n26756_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:579:46  */
  assign n26759_o = n26312_o[98];
  /* ../../HW/src/dp/dp_gen.vhd:579:66  */
  assign n26761_o = n26759_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:578:90  */
  assign n26762_o = n26761_o & n26758_o;
  /* ../../HW/src/dp/dp_gen.vhd:580:46  */
  assign n26763_o = n26312_o[196];
  /* ../../HW/src/dp/dp_gen.vhd:580:66  */
  assign n26765_o = n26763_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:579:90  */
  assign n26766_o = n26765_o & n26762_o;
  /* ../../HW/src/dp/dp_gen.vhd:581:46  */
  assign n26767_o = n26312_o[294];
  /* ../../HW/src/dp/dp_gen.vhd:581:66  */
  assign n26769_o = n26767_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:580:90  */
  assign n26770_o = n26769_o & n26766_o;
  /* ../../HW/src/dp/dp_gen.vhd:582:46  */
  assign n26771_o = n26312_o[392];
  /* ../../HW/src/dp/dp_gen.vhd:582:66  */
  assign n26773_o = n26771_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:581:90  */
  assign n26774_o = n26773_o & n26770_o;
  /* ../../HW/src/dp/dp_gen.vhd:583:39  */
  assign n26775_o = n26312_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:583:50  */
  assign n26777_o = n26775_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:582:90  */
  assign n26778_o = n26777_o & n26774_o;
  /* ../../HW/src/dp/dp_gen.vhd:584:44  */
  assign n26779_o = n26312_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:584:64  */
  assign n26781_o = n26779_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:583:111  */
  assign n26782_o = n26781_o & n26778_o;
  /* ../../HW/src/dp/dp_gen.vhd:585:48  */
  assign n26783_o = n26312_o[490];
  /* ../../HW/src/dp/dp_gen.vhd:585:68  */
  assign n26785_o = n26783_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:584:99  */
  assign n26786_o = n26785_o & n26782_o;
  /* ../../HW/src/dp/dp_gen.vhd:586:42  */
  assign n26787_o = n26312_o[593];
  /* ../../HW/src/dp/dp_gen.vhd:586:62  */
  assign n26789_o = n26787_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:585:103  */
  assign n26790_o = n26789_o & n26786_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:111  */
  assign n26791_o = n26755_o | n26790_o;
  /* ../../HW/src/dp/dp_gen.vhd:577:7  */
  assign n26794_o = n26791_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:569:7  */
  assign n26795_o = n26738_o ? n26752_o : n26794_o;
  /* ../../HW/src/dp/dp_gen.vhd:593:41  */
  assign n26797_o = pre_instruction_bus_id_dest_in == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:594:38  */
  assign n26798_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:594:49  */
  assign n26800_o = n26798_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:595:38  */
  assign n26801_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:595:49  */
  assign n26803_o = n26801_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:596:43  */
  assign n26804_o = n26313_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:596:63  */
  assign n26806_o = n26804_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:595:108  */
  assign n26807_o = n26806_o & n26803_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:108  */
  assign n26808_o = n26800_o | n26807_o;
  /* ../../HW/src/dp/dp_gen.vhd:594:11  */
  assign n26811_o = n26808_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:601:35  */
  assign n26812_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:601:46  */
  assign n26814_o = n26812_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:602:42  */
  assign n26815_o = n26313_o[0];
  /* ../../HW/src/dp/dp_gen.vhd:602:62  */
  assign n26817_o = n26815_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:603:42  */
  assign n26818_o = n26313_o[98];
  /* ../../HW/src/dp/dp_gen.vhd:603:62  */
  assign n26820_o = n26818_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:602:86  */
  assign n26821_o = n26820_o & n26817_o;
  /* ../../HW/src/dp/dp_gen.vhd:604:42  */
  assign n26822_o = n26313_o[196];
  /* ../../HW/src/dp/dp_gen.vhd:604:62  */
  assign n26824_o = n26822_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:603:86  */
  assign n26825_o = n26824_o & n26821_o;
  /* ../../HW/src/dp/dp_gen.vhd:605:42  */
  assign n26826_o = n26313_o[294];
  /* ../../HW/src/dp/dp_gen.vhd:605:62  */
  assign n26828_o = n26826_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:604:86  */
  assign n26829_o = n26828_o & n26825_o;
  /* ../../HW/src/dp/dp_gen.vhd:606:42  */
  assign n26830_o = n26313_o[392];
  /* ../../HW/src/dp/dp_gen.vhd:606:62  */
  assign n26832_o = n26830_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:605:86  */
  assign n26833_o = n26832_o & n26829_o;
  /* ../../HW/src/dp/dp_gen.vhd:607:35  */
  assign n26834_o = n26313_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:607:46  */
  assign n26836_o = n26834_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:606:86  */
  assign n26837_o = n26836_o & n26833_o;
  /* ../../HW/src/dp/dp_gen.vhd:608:40  */
  assign n26838_o = n26313_o[625];
  /* ../../HW/src/dp/dp_gen.vhd:608:60  */
  assign n26840_o = n26838_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:607:105  */
  assign n26841_o = n26840_o & n26837_o;
  /* ../../HW/src/dp/dp_gen.vhd:609:44  */
  assign n26842_o = n26313_o[490];
  /* ../../HW/src/dp/dp_gen.vhd:609:64  */
  assign n26844_o = n26842_o == 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:608:95  */
  assign n26845_o = n26844_o & n26841_o;
  /* ../../HW/src/dp/dp_gen.vhd:610:38  */
  assign n26846_o = n26313_o[593];
  /* ../../HW/src/dp/dp_gen.vhd:610:58  */
  assign n26848_o = n26846_o == 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:609:99  */
  assign n26849_o = n26848_o & n26845_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:105  */
  assign n26850_o = n26814_o | n26849_o;
  /* ../../HW/src/dp/dp_gen.vhd:601:5  */
  assign n26853_o = n26850_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:593:8  */
  assign n26854_o = n26797_o ? n26811_o : n26853_o;
  assign n26855_o = {n26795_o, n26643_o, n26491_o};
  assign n26857_o = {n26854_o, n26702_o, n26550_o};
  assign n26859_o = {n26719_o, n26567_o, n26415_o};
  assign n26861_o = {n26736_o, n26584_o, n26432_o};
  /* ../../HW/src/dp/dp_gen.vhd:627:21  */
  assign n26880_o = src_is_vector_r[0];
  /* ../../HW/src/dp/dp_gen.vhd:627:48  */
  assign n26881_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:627:51  */
  assign n26883_o = n26881_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:627:29  */
  assign n26884_o = n26880_o | n26883_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:95  */
  assign n26885_o = n26310_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:627:111  */
  assign n26886_o = ~n26885_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:69  */
  assign n26887_o = n26886_o & n26884_o;
  /* ../../HW/src/dp/dp_gen.vhd:628:21  */
  assign n26888_o = dst_is_vector_r[0];
  /* ../../HW/src/dp/dp_gen.vhd:628:48  */
  assign n26889_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:628:51  */
  assign n26891_o = n26889_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:628:29  */
  assign n26892_o = n26888_o | n26891_o;
  /* ../../HW/src/dp/dp_gen.vhd:628:93  */
  assign n26893_o = n26311_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:628:109  */
  assign n26894_o = ~n26893_o;
  /* ../../HW/src/dp/dp_gen.vhd:628:69  */
  assign n26895_o = n26894_o & n26892_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:117  */
  assign n26896_o = n26895_o & n26887_o;
  /* ../../HW/src/dp/dp_gen.vhd:631:35  */
  assign n26897_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:632:35  */
  assign n26898_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:633:23  */
  assign n26899_o = src_is_vector_r[1];
  /* ../../HW/src/dp/dp_gen.vhd:633:50  */
  assign n26900_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:633:53  */
  assign n26902_o = n26900_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:633:31  */
  assign n26903_o = n26899_o | n26902_o;
  /* ../../HW/src/dp/dp_gen.vhd:634:23  */
  assign n26904_o = dst_is_vector_r[1];
  /* ../../HW/src/dp/dp_gen.vhd:634:50  */
  assign n26905_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:634:53  */
  assign n26907_o = n26905_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:634:31  */
  assign n26908_o = n26904_o | n26907_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:71  */
  assign n26909_o = n26908_o & n26903_o;
  /* ../../HW/src/dp/dp_gen.vhd:637:35  */
  assign n26910_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:638:35  */
  assign n26911_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:639:23  */
  assign n26912_o = src_is_vector_r[2];
  /* ../../HW/src/dp/dp_gen.vhd:639:50  */
  assign n26913_o = src_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:639:53  */
  assign n26915_o = n26913_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:639:31  */
  assign n26916_o = n26912_o | n26915_o;
  /* ../../HW/src/dp/dp_gen.vhd:640:23  */
  assign n26917_o = dst_is_vector_r[2];
  /* ../../HW/src/dp/dp_gen.vhd:640:50  */
  assign n26918_o = dst_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:640:53  */
  assign n26920_o = n26918_o != 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:640:31  */
  assign n26921_o = n26917_o | n26920_o;
  /* ../../HW/src/dp/dp_gen.vhd:639:71  */
  assign n26922_o = n26921_o & n26916_o;
  /* ../../HW/src/dp/dp_gen.vhd:643:35  */
  assign n26923_o = src_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:644:35  */
  assign n26924_o = dst_is_scatter_r[5:4];
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n26927_o = n26922_o ? 3'b001 : 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n26930_o = n26922_o ? 3'b001 : 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n26932_o = n26922_o ? n26923_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:639:1  */
  assign n26934_o = n26922_o ? n26924_o : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n26936_o = n26909_o ? 3'b011 : n26927_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n26938_o = n26909_o ? 3'b011 : n26930_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n26939_o = n26909_o ? n26910_o : n26932_o;
  /* ../../HW/src/dp/dp_gen.vhd:633:1  */
  assign n26940_o = n26909_o ? n26911_o : n26934_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n26942_o = n26896_o ? 3'b111 : n26936_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n26944_o = n26896_o ? 3'b111 : n26938_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n26945_o = n26896_o ? n26897_o : n26939_o;
  /* ../../HW/src/dp/dp_gen.vhd:627:1  */
  assign n26946_o = n26896_o ? n26898_o : n26940_o;
  /* ../../HW/src/dp/dp_gen.vhd:658:31  */
  assign n26949_o = s_burstlen_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:659:56  */
  assign n26950_o = s_template_r[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:659:31  */
  assign n26951_o = s_burstpos_r + n26950_o;
  /* ../../HW/src/dp/dp_gen.vhd:660:40  */
  assign n26952_o = s_template_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:660:19  */
  assign n26953_o = s_i0_r + n26952_o;
  /* ../../HW/src/dp/dp_gen.vhd:661:40  */
  assign n26954_o = s_template_r[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:661:19  */
  assign n26955_o = s_i1_r + n26954_o;
  /* ../../HW/src/dp/dp_gen.vhd:662:40  */
  assign n26956_o = s_template_r[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:662:19  */
  assign n26957_o = s_i2_r + n26956_o;
  /* ../../HW/src/dp/dp_gen.vhd:663:40  */
  assign n26958_o = s_template_r[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:663:19  */
  assign n26959_o = s_i3_r + n26958_o;
  /* ../../HW/src/dp/dp_gen.vhd:664:40  */
  assign n26960_o = s_template_r[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:664:19  */
  assign n26961_o = s_i4_r + n26960_o;
  /* ../../HW/src/dp/dp_gen.vhd:666:57  */
  assign n26963_o = {1'b0, s_burstpos_stride_r};
  /* ../../HW/src/dp/dp_gen.vhd:666:43  */
  assign n26964_o = s_burstpos_start_r + n26963_o;
  /* ../../HW/src/dp/dp_gen.vhd:667:84  */
  assign n26965_o = s_template_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:667:45  */
  assign n26967_o = {1'b0, n26965_o};
  /* ../../HW/src/dp/dp_gen.vhd:667:31  */
  assign n26968_o = s_i0_start_r + n26967_o;
  /* ../../HW/src/dp/dp_gen.vhd:668:84  */
  assign n26969_o = s_template_r[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:668:45  */
  assign n26971_o = {1'b0, n26969_o};
  /* ../../HW/src/dp/dp_gen.vhd:668:31  */
  assign n26972_o = s_i1_start_r + n26971_o;
  /* ../../HW/src/dp/dp_gen.vhd:669:84  */
  assign n26973_o = s_template_r[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:669:45  */
  assign n26975_o = {1'b0, n26973_o};
  /* ../../HW/src/dp/dp_gen.vhd:669:31  */
  assign n26976_o = s_i2_start_r + n26975_o;
  /* ../../HW/src/dp/dp_gen.vhd:670:84  */
  assign n26977_o = s_template_r[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:670:45  */
  assign n26979_o = {1'b0, n26977_o};
  /* ../../HW/src/dp/dp_gen.vhd:670:31  */
  assign n26980_o = s_i3_start_r + n26979_o;
  /* ../../HW/src/dp/dp_gen.vhd:671:84  */
  assign n26981_o = s_template_r[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:671:45  */
  assign n26983_o = {1'b0, n26981_o};
  /* ../../HW/src/dp/dp_gen.vhd:671:31  */
  assign n26984_o = s_i4_start_r + n26983_o;
  /* ../../HW/src/dp/dp_gen.vhd:673:31  */
  assign n26986_o = s_i0_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:674:31  */
  assign n26988_o = s_i1_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:675:31  */
  assign n26990_o = s_i2_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:676:31  */
  assign n26992_o = s_i3_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:677:31  */
  assign n26994_o = s_i4_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:679:31  */
  assign n26996_o = d_burstlen_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:680:45  */
  assign n26997_o = d_template_r[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:680:31  */
  assign n26998_o = d_burstpos_r + n26997_o;
  /* ../../HW/src/dp/dp_gen.vhd:681:33  */
  assign n26999_o = d_template_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:681:19  */
  assign n27000_o = d_i0_r + n26999_o;
  /* ../../HW/src/dp/dp_gen.vhd:682:33  */
  assign n27001_o = d_template_r[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:682:19  */
  assign n27002_o = d_i1_r + n27001_o;
  /* ../../HW/src/dp/dp_gen.vhd:683:33  */
  assign n27003_o = d_template_r[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:683:19  */
  assign n27004_o = d_i2_r + n27003_o;
  /* ../../HW/src/dp/dp_gen.vhd:684:33  */
  assign n27005_o = d_template_r[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:684:19  */
  assign n27006_o = d_i3_r + n27005_o;
  /* ../../HW/src/dp/dp_gen.vhd:685:33  */
  assign n27007_o = d_template_r[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:685:19  */
  assign n27008_o = d_i4_r + n27007_o;
  /* ../../HW/src/dp/dp_gen.vhd:687:68  */
  assign n27009_o = d_template_r[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:687:97  */
  assign n27011_o = {n27009_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:687:20  */
  assign n27012_o = d_i0_r + n27011_o;
  /* ../../HW/src/dp/dp_gen.vhd:688:68  */
  assign n27013_o = d_template_r[120:98];
  /* ../../HW/src/dp/dp_gen.vhd:688:97  */
  assign n27015_o = {n27013_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:688:20  */
  assign n27016_o = d_i1_r + n27015_o;
  /* ../../HW/src/dp/dp_gen.vhd:689:68  */
  assign n27017_o = d_template_r[218:196];
  /* ../../HW/src/dp/dp_gen.vhd:689:97  */
  assign n27019_o = {n27017_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:689:20  */
  assign n27020_o = d_i2_r + n27019_o;
  /* ../../HW/src/dp/dp_gen.vhd:690:68  */
  assign n27021_o = d_template_r[316:294];
  /* ../../HW/src/dp/dp_gen.vhd:690:97  */
  assign n27023_o = {n27021_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:690:20  */
  assign n27024_o = d_i3_r + n27023_o;
  /* ../../HW/src/dp/dp_gen.vhd:691:68  */
  assign n27025_o = d_template_r[414:392];
  /* ../../HW/src/dp/dp_gen.vhd:691:97  */
  assign n27027_o = {n27025_o, 1'b0};
  /* ../../HW/src/dp/dp_gen.vhd:691:20  */
  assign n27028_o = d_i4_r + n27027_o;
  /* ../../HW/src/dp/dp_gen.vhd:693:31  */
  assign n27030_o = d_i0_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:694:31  */
  assign n27032_o = d_i1_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:695:31  */
  assign n27034_o = d_i2_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:696:31  */
  assign n27036_o = d_i3_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:697:31  */
  assign n27038_o = d_i4_count_r + 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:712:67  */
  assign n27041_o = ~s_gen_burstlen_progress_r;
  /* ../../HW/src/dp/dp_gen.vhd:712:39  */
  assign n27042_o = eof_rrrr | n27041_o;
  /* ../../HW/src/dp/dp_gen.vhd:712:20  */
  assign n27043_o = n27042_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:719:33  */
  assign n27046_o = waitreq_in & gen_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:719:49  */
  assign n27048_o = n27046_o != 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:719:16  */
  assign n27049_o = n27048_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:725:82  */
  assign n27052_o = s_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:725:53  */
  assign n27053_o = s_burstlen_r == n27052_o;
  /* ../../HW/src/dp/dp_gen.vhd:725:24  */
  assign n27054_o = n27053_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:726:84  */
  assign n27057_o = s_template_r[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:726:47  */
  assign n27058_o = s_i0_count_r == n27057_o;
  /* ../../HW/src/dp/dp_gen.vhd:726:18  */
  assign n27059_o = n27058_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:727:84  */
  assign n27062_o = s_template_r[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:727:47  */
  assign n27063_o = s_i1_count_r == n27062_o;
  /* ../../HW/src/dp/dp_gen.vhd:727:18  */
  assign n27064_o = n27063_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:728:84  */
  assign n27067_o = s_template_r[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:728:47  */
  assign n27068_o = s_i2_count_r == n27067_o;
  /* ../../HW/src/dp/dp_gen.vhd:728:18  */
  assign n27069_o = n27068_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:729:84  */
  assign n27072_o = s_template_r[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:729:47  */
  assign n27073_o = s_i3_count_r == n27072_o;
  /* ../../HW/src/dp/dp_gen.vhd:729:18  */
  assign n27074_o = n27073_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:730:84  */
  assign n27077_o = s_template_r[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:730:47  */
  assign n27078_o = s_i4_count_r == n27077_o;
  /* ../../HW/src/dp/dp_gen.vhd:730:18  */
  assign n27079_o = n27078_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:732:78  */
  assign n27082_o = s_template_r[71:48];
  /* ../../HW/src/dp/dp_gen.vhd:732:42  */
  assign n27083_o = $unsigned(s_i0_r) <= $unsigned(n27082_o);
  /* ../../HW/src/dp/dp_gen.vhd:732:136  */
  assign n27084_o = s_template_r[72];
  /* ../../HW/src/dp/dp_gen.vhd:732:153  */
  assign n27085_o = ~n27084_o;
  /* ../../HW/src/dp/dp_gen.vhd:732:108  */
  assign n27086_o = n27085_o & n27083_o;
  /* ../../HW/src/dp/dp_gen.vhd:732:19  */
  assign n27087_o = n27086_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:733:78  */
  assign n27090_o = s_template_r[169:146];
  /* ../../HW/src/dp/dp_gen.vhd:733:42  */
  assign n27091_o = $unsigned(s_i1_r) <= $unsigned(n27090_o);
  /* ../../HW/src/dp/dp_gen.vhd:733:136  */
  assign n27092_o = s_template_r[170];
  /* ../../HW/src/dp/dp_gen.vhd:733:153  */
  assign n27093_o = ~n27092_o;
  /* ../../HW/src/dp/dp_gen.vhd:733:108  */
  assign n27094_o = n27093_o & n27091_o;
  /* ../../HW/src/dp/dp_gen.vhd:733:19  */
  assign n27095_o = n27094_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:734:78  */
  assign n27098_o = s_template_r[267:244];
  /* ../../HW/src/dp/dp_gen.vhd:734:42  */
  assign n27099_o = $unsigned(s_i2_r) <= $unsigned(n27098_o);
  /* ../../HW/src/dp/dp_gen.vhd:734:136  */
  assign n27100_o = s_template_r[268];
  /* ../../HW/src/dp/dp_gen.vhd:734:153  */
  assign n27101_o = ~n27100_o;
  /* ../../HW/src/dp/dp_gen.vhd:734:108  */
  assign n27102_o = n27101_o & n27099_o;
  /* ../../HW/src/dp/dp_gen.vhd:734:19  */
  assign n27103_o = n27102_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:735:78  */
  assign n27106_o = s_template_r[365:342];
  /* ../../HW/src/dp/dp_gen.vhd:735:42  */
  assign n27107_o = $unsigned(s_i3_r) <= $unsigned(n27106_o);
  /* ../../HW/src/dp/dp_gen.vhd:735:136  */
  assign n27108_o = s_template_r[366];
  /* ../../HW/src/dp/dp_gen.vhd:735:153  */
  assign n27109_o = ~n27108_o;
  /* ../../HW/src/dp/dp_gen.vhd:735:108  */
  assign n27110_o = n27109_o & n27107_o;
  /* ../../HW/src/dp/dp_gen.vhd:735:19  */
  assign n27111_o = n27110_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:736:78  */
  assign n27114_o = s_template_r[463:440];
  /* ../../HW/src/dp/dp_gen.vhd:736:42  */
  assign n27115_o = $unsigned(s_i4_r) <= $unsigned(n27114_o);
  /* ../../HW/src/dp/dp_gen.vhd:736:136  */
  assign n27116_o = s_template_r[464];
  /* ../../HW/src/dp/dp_gen.vhd:736:153  */
  assign n27117_o = ~n27116_o;
  /* ../../HW/src/dp/dp_gen.vhd:736:108  */
  assign n27118_o = n27117_o & n27115_o;
  /* ../../HW/src/dp/dp_gen.vhd:736:19  */
  assign n27119_o = n27118_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:737:85  */
  assign n27122_o = s_template_r[513:490];
  /* ../../HW/src/dp/dp_gen.vhd:737:51  */
  assign n27123_o = $unsigned(s_burstpos_r) <= $unsigned(n27122_o);
  /* ../../HW/src/dp/dp_gen.vhd:737:141  */
  assign n27124_o = s_template_r[514];
  /* ../../HW/src/dp/dp_gen.vhd:737:158  */
  assign n27125_o = ~n27124_o;
  /* ../../HW/src/dp/dp_gen.vhd:737:115  */
  assign n27126_o = n27125_o & n27123_o;
  /* ../../HW/src/dp/dp_gen.vhd:737:22  */
  assign n27127_o = n27126_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:739:37  */
  assign n27129_o = s_i0_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:739:21  */
  assign n27130_o = ~n27129_o;
  /* ../../HW/src/dp/dp_gen.vhd:740:37  */
  assign n27131_o = s_i1_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:740:21  */
  assign n27132_o = ~n27131_o;
  /* ../../HW/src/dp/dp_gen.vhd:741:37  */
  assign n27133_o = s_i2_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:741:21  */
  assign n27134_o = ~n27133_o;
  /* ../../HW/src/dp/dp_gen.vhd:742:37  */
  assign n27135_o = s_i3_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:742:21  */
  assign n27136_o = ~n27135_o;
  /* ../../HW/src/dp/dp_gen.vhd:743:37  */
  assign n27137_o = s_i4_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:743:21  */
  assign n27138_o = ~n27137_o;
  /* ../../HW/src/dp/dp_gen.vhd:744:61  */
  assign n27140_o = {{1{s_burstpos_stride_r[23]}}, s_burstpos_stride_r}; // sext
  /* ../../HW/src/dp/dp_gen.vhd:744:61  */
  assign n27141_o = s_burstpos_start_r + n27140_o;
  /* ../../HW/src/dp/dp_gen.vhd:744:91  */
  assign n27143_o = $signed(n27141_o) >= $signed(25'b0000000000000000000000001);
  /* ../../HW/src/dp/dp_gen.vhd:744:28  */
  assign n27144_o = n27143_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:746:77  */
  assign n27147_o = d_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:746:53  */
  assign n27148_o = d_burstlen_r == n27147_o;
  /* ../../HW/src/dp/dp_gen.vhd:746:24  */
  assign n27149_o = n27148_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:747:71  */
  assign n27152_o = d_template_r[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:747:47  */
  assign n27153_o = d_i0_count_r == n27152_o;
  /* ../../HW/src/dp/dp_gen.vhd:747:18  */
  assign n27154_o = n27153_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:748:71  */
  assign n27157_o = d_template_r[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:748:47  */
  assign n27158_o = d_i1_count_r == n27157_o;
  /* ../../HW/src/dp/dp_gen.vhd:748:18  */
  assign n27159_o = n27158_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:749:71  */
  assign n27162_o = d_template_r[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:749:47  */
  assign n27163_o = d_i2_count_r == n27162_o;
  /* ../../HW/src/dp/dp_gen.vhd:749:18  */
  assign n27164_o = n27163_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:750:71  */
  assign n27167_o = d_template_r[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:750:47  */
  assign n27168_o = d_i3_count_r == n27167_o;
  /* ../../HW/src/dp/dp_gen.vhd:750:18  */
  assign n27169_o = n27168_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:751:71  */
  assign n27172_o = d_template_r[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:751:47  */
  assign n27173_o = d_i4_count_r == n27172_o;
  /* ../../HW/src/dp/dp_gen.vhd:751:18  */
  assign n27174_o = n27173_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:753:78  */
  assign n27177_o = d_template_r[71:48];
  /* ../../HW/src/dp/dp_gen.vhd:753:42  */
  assign n27178_o = $unsigned(d_i0_r) <= $unsigned(n27177_o);
  /* ../../HW/src/dp/dp_gen.vhd:753:136  */
  assign n27179_o = d_template_r[72];
  /* ../../HW/src/dp/dp_gen.vhd:753:153  */
  assign n27180_o = ~n27179_o;
  /* ../../HW/src/dp/dp_gen.vhd:753:108  */
  assign n27181_o = n27180_o & n27178_o;
  /* ../../HW/src/dp/dp_gen.vhd:753:19  */
  assign n27182_o = n27181_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:754:78  */
  assign n27185_o = d_template_r[169:146];
  /* ../../HW/src/dp/dp_gen.vhd:754:42  */
  assign n27186_o = $unsigned(d_i1_r) <= $unsigned(n27185_o);
  /* ../../HW/src/dp/dp_gen.vhd:754:136  */
  assign n27187_o = d_template_r[170];
  /* ../../HW/src/dp/dp_gen.vhd:754:153  */
  assign n27188_o = ~n27187_o;
  /* ../../HW/src/dp/dp_gen.vhd:754:108  */
  assign n27189_o = n27188_o & n27186_o;
  /* ../../HW/src/dp/dp_gen.vhd:754:19  */
  assign n27190_o = n27189_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:755:78  */
  assign n27193_o = d_template_r[267:244];
  /* ../../HW/src/dp/dp_gen.vhd:755:42  */
  assign n27194_o = $unsigned(d_i2_r) <= $unsigned(n27193_o);
  /* ../../HW/src/dp/dp_gen.vhd:755:136  */
  assign n27195_o = d_template_r[268];
  /* ../../HW/src/dp/dp_gen.vhd:755:153  */
  assign n27196_o = ~n27195_o;
  /* ../../HW/src/dp/dp_gen.vhd:755:108  */
  assign n27197_o = n27196_o & n27194_o;
  /* ../../HW/src/dp/dp_gen.vhd:755:19  */
  assign n27198_o = n27197_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:756:78  */
  assign n27201_o = d_template_r[365:342];
  /* ../../HW/src/dp/dp_gen.vhd:756:42  */
  assign n27202_o = $unsigned(d_i3_r) <= $unsigned(n27201_o);
  /* ../../HW/src/dp/dp_gen.vhd:756:136  */
  assign n27203_o = d_template_r[366];
  /* ../../HW/src/dp/dp_gen.vhd:756:153  */
  assign n27204_o = ~n27203_o;
  /* ../../HW/src/dp/dp_gen.vhd:756:108  */
  assign n27205_o = n27204_o & n27202_o;
  /* ../../HW/src/dp/dp_gen.vhd:756:19  */
  assign n27206_o = n27205_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:757:78  */
  assign n27209_o = d_template_r[463:440];
  /* ../../HW/src/dp/dp_gen.vhd:757:42  */
  assign n27210_o = $unsigned(d_i4_r) <= $unsigned(n27209_o);
  /* ../../HW/src/dp/dp_gen.vhd:757:136  */
  assign n27211_o = d_template_r[464];
  /* ../../HW/src/dp/dp_gen.vhd:757:153  */
  assign n27212_o = ~n27211_o;
  /* ../../HW/src/dp/dp_gen.vhd:757:108  */
  assign n27213_o = n27212_o & n27210_o;
  /* ../../HW/src/dp/dp_gen.vhd:757:19  */
  assign n27214_o = n27213_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:758:76  */
  assign n27217_o = d_burst_max_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:758:51  */
  assign n27218_o = $unsigned(d_burstpos_r) <= $unsigned(n27217_o);
  /* ../../HW/src/dp/dp_gen.vhd:758:123  */
  assign n27219_o = d_burst_max_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:758:140  */
  assign n27220_o = ~n27219_o;
  /* ../../HW/src/dp/dp_gen.vhd:758:106  */
  assign n27221_o = n27220_o & n27218_o;
  /* ../../HW/src/dp/dp_gen.vhd:758:22  */
  assign n27222_o = n27221_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:776:16  */
  assign n27234_o = ~reset_in;
  /* ../../HW/src/dp/dp_gen.vhd:915:24  */
  assign n27236_o = ~waitreq;
  /* ../../HW/src/dp/dp_gen.vhd:920:40  */
  assign n27238_o = dp_src_bus_id_rrr == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:920:20  */
  assign n27240_o = n27238_o ? running_rrr : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:920:40  */
  assign n27242_o = dp_src_bus_id_rrr == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:920:20  */
  assign n27244_o = n27242_o ? running_rrr : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:920:40  */
  assign n27246_o = dp_src_bus_id_rrr == 2'b10;
  /* ../../HW/src/dp/dp_gen.vhd:920:20  */
  assign n27248_o = n27246_o ? running_rrr : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:971:36  */
  assign n27252_o = s_i0_r + s_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:971:43  */
  assign n27253_o = n27252_o + s_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:972:52  */
  assign n27254_o = s_template_r[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:974:46  */
  assign n27255_o = s_template_r[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:975:48  */
  assign n27256_o = s_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:975:76  */
  assign n27257_o = n27256_o - s_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:976:42  */
  assign n27258_o = s_burstpos_r + s_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:976:49  */
  assign n27259_o = n27258_o + s_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:977:39  */
  assign n27260_o = s_temp1_r + s_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:979:27  */
  assign n27261_o = {8'b0, s_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:979:75  */
  assign n27262_o = n27261_o + s_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:981:43  */
  assign n27264_o = n27262_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:980:17  */
  assign n27265_o = src_double_rrr ? n27264_o : n27262_o;
  /* ../../HW/src/dp/dp_gen.vhd:985:37  */
  assign n27269_o = $unsigned(s_gen_burstlen_r) > $unsigned(n29586_o);
  /* ../../HW/src/dp/dp_gen.vhd:985:17  */
  assign n27273_o = n27269_o ? n29593_o : s_gen_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:991:34  */
  assign n27275_o = n27273_o == 5'b00000;
  /* ../../HW/src/dp/dp_gen.vhd:991:17  */
  assign n27278_o = n27275_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:1001:40  */
  assign n27279_o = {3'b0, s_burstpos_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1002:65  */
  assign n27280_o = s_burst_actual_max_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1002:38  */
  assign n27281_o = {3'b0, n27280_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1002:110  */
  assign n27282_o = n27281_o - n27279_o;
  /* ../../HW/src/dp/dp_gen.vhd:1002:122  */
  assign n27284_o = n27282_o + 27'b000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1004:39  */
  assign n27286_o = n27284_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1003:17  */
  assign n27287_o = src_double_r ? n27286_o : n27284_o;
  /* ../../HW/src/dp/dp_gen.vhd:1007:36  */
  assign n27288_o = s_burstpos_end_r[26];
  /* ../../HW/src/dp/dp_gen.vhd:1010:39  */
  assign n27289_o = s_burstpos_end_r[26:4];
  /* ../../HW/src/dp/dp_gen.vhd:1010:94  */
  assign n27291_o = n27289_o == 23'b00000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1012:57  */
  assign n27292_o = s_burstpos_end_r[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1010:17  */
  assign n27294_o = n27291_o ? n27292_o : 4'b1111;
  /* ../../HW/src/dp/dp_gen.vhd:1007:17  */
  assign n27296_o = n27288_o ? 4'b0000 : n27294_o;
  /* ../../HW/src/dp/dp_gen.vhd:1020:55  */
  assign n27297_o = s_bufsize_rr[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:1020:36  */
  assign n27298_o = {2'b0, n27297_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1020:111  */
  assign n27299_o = {1'b0, s_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1020:103  */
  assign n27300_o = n27298_o - n27299_o;
  /* ../../HW/src/dp/dp_gen.vhd:1022:41  */
  assign n27302_o = n27300_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1021:17  */
  assign n27303_o = src_double_rrr ? n27302_o : n27300_o;
  /* ../../HW/src/dp/dp_gen.vhd:1024:29  */
  assign n27305_o = $signed(n27303_o) <= $signed(25'b0000000000000000000000000);
  /* ../../HW/src/dp/dp_gen.vhd:1026:44  */
  assign n27306_o = {21'b0, s_burstpos_end_rr};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1026:42  */
  assign n27307_o = $unsigned(n27303_o) > $unsigned(n27306_o);
  /* ../../HW/src/dp/dp_gen.vhd:1029:59  */
  assign n27308_o = n27303_o[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1026:17  */
  assign n27309_o = n27307_o ? s_burstpos_end_rr : n27308_o;
  /* ../../HW/src/dp/dp_gen.vhd:1024:17  */
  assign n27311_o = n27305_o ? 4'b0000 : n27309_o;
  /* ../../HW/src/dp/dp_gen.vhd:1032:89  */
  assign n27313_o = s_template_r[512:490];
  /* ../../HW/src/dp/dp_gen.vhd:1032:47  */
  assign n27315_o = {1'b0, n27313_o};
  /* ../../HW/src/dp/dp_gen.vhd:1032:120  */
  assign n27316_o = n27315_o - s_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1033:42  */
  assign n27318_o = src_vector_r == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1034:106  */
  assign n27319_o = n27316_o[23:1];
  /* ../../HW/src/dp/dp_gen.vhd:1036:45  */
  assign n27322_o = src_vector_r == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1037:106  */
  assign n27323_o = n27316_o[23:2];
  /* ../../HW/src/dp/dp_gen.vhd:1039:45  */
  assign n27326_o = src_vector_r == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1040:104  */
  assign n27327_o = n27316_o[23:3];
  assign n27329_o = {3'b000, n27327_o};
  /* ../../HW/src/dp/dp_gen.vhd:1039:17  */
  assign n27330_o = n27326_o ? n27329_o : n27316_o;
  assign n27331_o = {2'b00, n27323_o};
  /* ../../HW/src/dp/dp_gen.vhd:1036:17  */
  assign n27332_o = n27322_o ? n27331_o : n27330_o;
  assign n27333_o = {1'b0, n27319_o};
  /* ../../HW/src/dp/dp_gen.vhd:1033:17  */
  assign n27334_o = n27318_o ? n27333_o : n27332_o;
  /* ../../HW/src/dp/dp_gen.vhd:1045:42  */
  assign n27335_o = s_i0_valid & s_i1_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:57  */
  assign n27336_o = n27335_o & s_i2_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:72  */
  assign n27337_o = n27336_o & s_i3_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:87  */
  assign n27338_o = n27337_o & s_i4_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:102  */
  assign n27339_o = n27338_o & s_burst_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:48  */
  assign n27340_o = s_i0_start_valid & s_i1_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:69  */
  assign n27341_o = n27340_o & s_i2_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:90  */
  assign n27342_o = n27341_o & s_i3_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:111  */
  assign n27343_o = n27342_o & s_i4_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1046:132  */
  assign n27344_o = n27343_o & s_burst_start_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1045:121  */
  assign n27345_o = n27339_o & n27344_o;
  /* ../../HW/src/dp/dp_gen.vhd:1047:29  */
  assign n27346_o = ~s_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:1049:45  */
  assign n27348_o = src_is_burst_rr & 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:1050:33  */
  assign n27349_o = s_temp3_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1050:78  */
  assign n27351_o = n27349_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1051:32  */
  assign n27352_o = s_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1051:62  */
  assign n27354_o = n27352_o != 5'b11111;
  /* ../../HW/src/dp/dp_gen.vhd:1050:129  */
  assign n27355_o = n27354_o & n27351_o;
  /* ../../HW/src/dp/dp_gen.vhd:1052:48  */
  assign n27356_o = s_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1050:20  */
  assign n27358_o = n27355_o ? n27356_o : 5'b11110;
  /* ../../HW/src/dp/dp_gen.vhd:1056:38  */
  assign n27359_o = s_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1058:41  */
  assign n27360_o = s_burstremain_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1058:92  */
  assign n27362_o = n27360_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1059:53  */
  assign n27363_o = s_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1059:36  */
  assign n27364_o = $unsigned(n27358_o) > $unsigned(n27363_o);
  /* ../../HW/src/dp/dp_gen.vhd:1058:149  */
  assign n27365_o = n27364_o & n27362_o;
  /* ../../HW/src/dp/dp_gen.vhd:1060:58  */
  assign n27366_o = s_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1060:88  */
  assign n27368_o = n27366_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1062:55  */
  assign n27370_o = n27358_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1058:20  */
  assign n27371_o = n27365_o ? n27368_o : n27370_o;
  /* ../../HW/src/dp/dp_gen.vhd:1056:20  */
  assign n27373_o = n27359_o ? 5'b00000 : n27371_o;
  /* ../../HW/src/dp/dp_gen.vhd:1065:38  */
  assign n27374_o = s_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1065:20  */
  assign n27377_o = n27374_o ? 5'b00000 : 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1049:17  */
  assign n27378_o = n27348_o ? n27373_o : n27377_o;
  /* ../../HW/src/dp/dp_gen.vhd:1047:17  */
  assign n27381_o = n27346_o ? 5'b00000 : n27378_o;
  /* ../../HW/src/dp/dp_gen.vhd:1103:84  */
  assign n27383_o = src_vector_rrr[1:0];
  assign n27385_o = {n27383_o, 1'b1};
  /* ../../HW/src/dp/dp_gen.vhd:1102:17  */
  assign n27386_o = src_double_rrr ? n27385_o : src_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:1112:38  */
  assign n27387_o = s_burstpos_start_r[24];
  /* ../../HW/src/dp/dp_gen.vhd:1112:67  */
  assign n27388_o = ~n27387_o;
  /* ../../HW/src/dp/dp_gen.vhd:1115:41  */
  assign n27389_o = s_burstpos_start_r[24:3];
  /* ../../HW/src/dp/dp_gen.vhd:1115:96  */
  assign n27391_o = n27389_o == 22'b1111111111111111111111;
  /* ../../HW/src/dp/dp_gen.vhd:1117:61  */
  assign n27392_o = s_burstpos_start_r[3:0];
  assign n27395_o = {1'b1, 3'b000};
  /* ../../HW/src/dp/dp_gen.vhd:1115:17  */
  assign n27396_o = n27391_o ? n27392_o : n27395_o;
  /* ../../HW/src/dp/dp_gen.vhd:1112:17  */
  assign n27398_o = n27388_o ? 4'b0000 : n27396_o;
  /* ../../HW/src/dp/dp_gen.vhd:1129:84  */
  assign n27399_o = dst_vector_rrr[1:0];
  assign n27401_o = {n27399_o, 1'b1};
  /* ../../HW/src/dp/dp_gen.vhd:1128:17  */
  assign n27402_o = dst_double_rrr ? n27401_o : dst_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:1155:52  */
  assign n27403_o = d_template_r[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:1157:36  */
  assign n27404_o = d_i0_r + d_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:1157:43  */
  assign n27405_o = n27404_o + d_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:1158:43  */
  assign n27406_o = d_template_r[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:1159:43  */
  assign n27407_o = d_template_r[648:625];
  /* ../../HW/src/dp/dp_gen.vhd:1159:48  */
  assign n27408_o = n27407_o - d_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1160:42  */
  assign n27409_o = d_burstpos_r + d_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:1160:49  */
  assign n27410_o = n27409_o + d_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1161:39  */
  assign n27411_o = d_temp1_r + d_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1164:27  */
  assign n27412_o = {8'b0, d_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1164:75  */
  assign n27413_o = n27412_o + d_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:1166:43  */
  assign n27415_o = n27413_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1165:17  */
  assign n27416_o = dst_double_rrr ? n27415_o : n27413_o;
  /* ../../HW/src/dp/dp_gen.vhd:1173:40  */
  assign n27417_o = {3'b0, d_burstpos_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1174:58  */
  assign n27418_o = d_burst_max_r[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1174:38  */
  assign n27419_o = {3'b0, n27418_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1174:103  */
  assign n27420_o = n27419_o - n27417_o;
  /* ../../HW/src/dp/dp_gen.vhd:1174:115  */
  assign n27422_o = n27420_o + 27'b000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1176:39  */
  assign n27424_o = n27422_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1175:17  */
  assign n27425_o = dst_double_r ? n27424_o : n27422_o;
  /* ../../HW/src/dp/dp_gen.vhd:1179:36  */
  assign n27426_o = d_burstpos_end_r[26];
  /* ../../HW/src/dp/dp_gen.vhd:1181:39  */
  assign n27427_o = d_burstpos_end_r[26:4];
  /* ../../HW/src/dp/dp_gen.vhd:1181:94  */
  assign n27429_o = n27427_o == 23'b00000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1182:57  */
  assign n27430_o = d_burstpos_end_r[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1181:17  */
  assign n27432_o = n27429_o ? n27430_o : 4'b1111;
  /* ../../HW/src/dp/dp_gen.vhd:1179:17  */
  assign n27434_o = n27426_o ? 4'b0000 : n27432_o;
  /* ../../HW/src/dp/dp_gen.vhd:1188:55  */
  assign n27435_o = d_bufsize_rr[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:1188:36  */
  assign n27436_o = {2'b0, n27435_o};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1188:111  */
  assign n27437_o = {1'b0, d_temp5_r};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1188:103  */
  assign n27438_o = n27436_o - n27437_o;
  /* ../../HW/src/dp/dp_gen.vhd:1190:41  */
  assign n27440_o = n27438_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1189:17  */
  assign n27441_o = dst_double_rrr ? n27440_o : n27438_o;
  /* ../../HW/src/dp/dp_gen.vhd:1192:29  */
  assign n27443_o = $signed(n27441_o) <= $signed(25'b0000000000000000000000000);
  /* ../../HW/src/dp/dp_gen.vhd:1194:44  */
  assign n27444_o = {21'b0, d_burstpos_end_rr};  //  uext
  /* ../../HW/src/dp/dp_gen.vhd:1194:42  */
  assign n27445_o = $unsigned(n27441_o) > $unsigned(n27444_o);
  /* ../../HW/src/dp/dp_gen.vhd:1197:59  */
  assign n27446_o = n27441_o[3:0];
  /* ../../HW/src/dp/dp_gen.vhd:1194:17  */
  assign n27447_o = n27445_o ? d_burstpos_end_rr : n27446_o;
  /* ../../HW/src/dp/dp_gen.vhd:1192:17  */
  assign n27449_o = n27443_o ? 4'b0000 : n27447_o;
  /* ../../HW/src/dp/dp_gen.vhd:1201:79  */
  assign n27451_o = d_burst_max_r[22:0];
  /* ../../HW/src/dp/dp_gen.vhd:1201:47  */
  assign n27453_o = {1'b0, n27451_o};
  /* ../../HW/src/dp/dp_gen.vhd:1201:109  */
  assign n27454_o = n27453_o - d_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1202:42  */
  assign n27456_o = dst_vector_r == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1203:106  */
  assign n27457_o = n27454_o[23:1];
  /* ../../HW/src/dp/dp_gen.vhd:1205:45  */
  assign n27460_o = dst_vector_r == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1206:106  */
  assign n27461_o = n27454_o[23:2];
  /* ../../HW/src/dp/dp_gen.vhd:1208:45  */
  assign n27464_o = dst_vector_r == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1209:104  */
  assign n27465_o = n27454_o[23:3];
  assign n27467_o = {3'b000, n27465_o};
  /* ../../HW/src/dp/dp_gen.vhd:1208:17  */
  assign n27468_o = n27464_o ? n27467_o : n27454_o;
  assign n27469_o = {2'b00, n27461_o};
  /* ../../HW/src/dp/dp_gen.vhd:1205:17  */
  assign n27470_o = n27460_o ? n27469_o : n27468_o;
  assign n27471_o = {1'b0, n27457_o};
  /* ../../HW/src/dp/dp_gen.vhd:1202:17  */
  assign n27472_o = n27456_o ? n27471_o : n27470_o;
  /* ../../HW/src/dp/dp_gen.vhd:1214:42  */
  assign n27473_o = d_i0_valid & d_i1_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:57  */
  assign n27474_o = n27473_o & d_i2_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:72  */
  assign n27475_o = n27474_o & d_i3_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:87  */
  assign n27476_o = n27475_o & d_i4_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1214:102  */
  assign n27477_o = n27476_o & d_burst_valid;
  /* ../../HW/src/dp/dp_gen.vhd:1215:29  */
  assign n27478_o = ~d_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:1217:43  */
  assign n27480_o = dst_is_burst_rr & 1'b1;
  /* ../../HW/src/dp/dp_gen.vhd:1218:34  */
  assign n27481_o = d_temp3_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1218:79  */
  assign n27483_o = n27481_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1219:34  */
  assign n27484_o = d_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1219:64  */
  assign n27486_o = n27484_o != 5'b11111;
  /* ../../HW/src/dp/dp_gen.vhd:1218:130  */
  assign n27487_o = n27486_o & n27483_o;
  /* ../../HW/src/dp/dp_gen.vhd:1220:50  */
  assign n27488_o = d_temp3_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1218:21  */
  assign n27490_o = n27487_o ? n27488_o : 5'b11110;
  /* ../../HW/src/dp/dp_gen.vhd:1224:39  */
  assign n27491_o = d_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1226:42  */
  assign n27492_o = d_burstremain_r[23:5];
  /* ../../HW/src/dp/dp_gen.vhd:1226:93  */
  assign n27494_o = n27492_o == 19'b0000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1227:57  */
  assign n27495_o = d_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1227:40  */
  assign n27496_o = $unsigned(n27490_o) > $unsigned(n27495_o);
  /* ../../HW/src/dp/dp_gen.vhd:1226:150  */
  assign n27497_o = n27496_o & n27494_o;
  /* ../../HW/src/dp/dp_gen.vhd:1228:60  */
  assign n27498_o = d_burstremain_r[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:1228:90  */
  assign n27500_o = n27498_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1230:57  */
  assign n27502_o = n27490_o + 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1226:21  */
  assign n27503_o = n27497_o ? n27500_o : n27502_o;
  /* ../../HW/src/dp/dp_gen.vhd:1224:21  */
  assign n27505_o = n27491_o ? 5'b00000 : n27503_o;
  /* ../../HW/src/dp/dp_gen.vhd:1233:39  */
  assign n27506_o = d_burstremain_r[23];
  /* ../../HW/src/dp/dp_gen.vhd:1233:21  */
  assign n27509_o = n27506_o ? 5'b00000 : 5'b00001;
  /* ../../HW/src/dp/dp_gen.vhd:1217:17  */
  assign n27510_o = n27480_o ? n27505_o : n27509_o;
  /* ../../HW/src/dp/dp_gen.vhd:1215:17  */
  assign n27513_o = n27478_o ? 5'b00000 : n27510_o;
  assign n27536_o = {n27248_o, n27244_o, n27240_o};
  /* ../../HW/src/dp/dp_gen.vhd:915:14  */
  assign n27632_o = n27236_o ? n29579_o : n29600_o;
  /* ../../HW/src/dp/dp_gen.vhd:1252:10  */
  always @*
    n28032_burst_min_v = n29128_q; // (isignal)
  initial
    n28032_burst_min_v = 25'bX;
  /* ../../HW/src/dp/dp_gen.vhd:1256:16  */
  assign n28038_o = ~reset_in;
  /* ../../HW/src/dp/dp_gen.vhd:1333:21  */
  assign n28040_o = ~waitreq;
  /* ../../HW/src/dp/dp_gen.vhd:1333:42  */
  assign n28041_o = instruction_valid_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1333:27  */
  assign n28042_o = n28040_o | n28041_o;
  /* ../../HW/src/dp/dp_gen.vhd:1335:16  */
  assign n28046_o = instruction_valid_in ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1347:65  */
  assign n28047_o = n26310_o[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1348:71  */
  assign n28048_o = n26310_o[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:1349:69  */
  assign n28049_o = n26310_o[72:48];
  /* ../../HW/src/dp/dp_gen.vhd:1350:69  */
  assign n28050_o = n26310_o[97:73];
  /* ../../HW/src/dp/dp_gen.vhd:1351:65  */
  assign n28051_o = n26310_o[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:1352:71  */
  assign n28052_o = n26310_o[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:1353:69  */
  assign n28053_o = n26310_o[170:146];
  /* ../../HW/src/dp/dp_gen.vhd:1354:69  */
  assign n28054_o = n26310_o[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1355:65  */
  assign n28055_o = n26310_o[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:1356:71  */
  assign n28056_o = n26310_o[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:1357:69  */
  assign n28057_o = n26310_o[268:244];
  /* ../../HW/src/dp/dp_gen.vhd:1358:69  */
  assign n28058_o = n26310_o[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1359:65  */
  assign n28059_o = n26310_o[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:1360:71  */
  assign n28060_o = n26310_o[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:1361:69  */
  assign n28061_o = n26310_o[366:342];
  /* ../../HW/src/dp/dp_gen.vhd:1362:69  */
  assign n28062_o = n26310_o[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1363:65  */
  assign n28063_o = n26310_o[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:1364:71  */
  assign n28064_o = n26310_o[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:1365:69  */
  assign n28065_o = n26310_o[464:440];
  /* ../../HW/src/dp/dp_gen.vhd:1366:69  */
  assign n28066_o = n26310_o[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1367:135  */
  assign n28067_o = n26310_o[514:493];
  /* ../../HW/src/dp/dp_gen.vhd:1369:82  */
  assign n28068_o = n26310_o[490];
  /* ../../HW/src/dp/dp_gen.vhd:1369:99  */
  assign n28069_o = src_vector[0];
  /* ../../HW/src/dp/dp_gen.vhd:1369:86  */
  assign n28070_o = n28068_o | n28069_o;
  /* ../../HW/src/dp/dp_gen.vhd:1369:82  */
  assign n28071_o = n26310_o[491];
  /* ../../HW/src/dp/dp_gen.vhd:1369:99  */
  assign n28072_o = src_vector[1];
  /* ../../HW/src/dp/dp_gen.vhd:1369:86  */
  assign n28073_o = n28071_o | n28072_o;
  /* ../../HW/src/dp/dp_gen.vhd:1369:82  */
  assign n28074_o = n26310_o[492];
  /* ../../HW/src/dp/dp_gen.vhd:1369:99  */
  assign n28075_o = src_vector[2];
  /* ../../HW/src/dp/dp_gen.vhd:1369:86  */
  assign n28076_o = n28074_o | n28075_o;
  /* ../../HW/src/dp/dp_gen.vhd:1371:65  */
  assign n28077_o = n26310_o[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1373:65  */
  assign n28078_o = n26310_o[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:1374:61  */
  assign n28079_o = n26310_o[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:1375:71  */
  assign n28080_o = n26310_o[775:752];
  /* ../../HW/src/dp/dp_gen.vhd:1377:32  */
  assign n28082_o = src_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1378:128  */
  assign n28083_o = n26310_o[648:628];
  /* ../../HW/src/dp/dp_gen.vhd:1380:35  */
  assign n28086_o = src_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1381:130  */
  assign n28087_o = n26310_o[648:627];
  /* ../../HW/src/dp/dp_gen.vhd:1383:35  */
  assign n28090_o = src_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1384:130  */
  assign n28091_o = n26310_o[648:626];
  /* ../../HW/src/dp/dp_gen.vhd:1387:66  */
  assign n28093_o = n26310_o[648:625];
  assign n28094_o = {1'b0, n28091_o};
  /* ../../HW/src/dp/dp_gen.vhd:1383:19  */
  assign n28095_o = n28090_o ? n28094_o : n28093_o;
  assign n28096_o = {2'b00, n28087_o};
  /* ../../HW/src/dp/dp_gen.vhd:1380:19  */
  assign n28097_o = n28086_o ? n28096_o : n28095_o;
  assign n28098_o = {3'b000, n28083_o};
  /* ../../HW/src/dp/dp_gen.vhd:1377:19  */
  assign n28099_o = n28082_o ? n28098_o : n28097_o;
  /* ../../HW/src/dp/dp_gen.vhd:1391:59  */
  assign n28100_o = n26310_o[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1391:69  */
  assign n28102_o = n28100_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1393:59  */
  assign n28103_o = n26310_o[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1390:19  */
  assign n28104_o = source_double_precision ? n28102_o : n28103_o;
  /* ../../HW/src/dp/dp_gen.vhd:1397:44  */
  assign n28105_o = n26310_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1397:55  */
  assign n28107_o = n28105_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1397:19  */
  assign n28110_o = n28107_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1402:32  */
  assign n28112_o = src_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1403:41  */
  assign n28113_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1403:44  */
  assign n28115_o = n28113_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1405:44  */
  assign n28116_o = src_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1405:47  */
  assign n28118_o = n28116_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1405:22  */
  assign n28121_o = n28118_o ? 24'b000000000000000001000000 : 24'b000000000000100000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1403:22  */
  assign n28123_o = n28115_o ? 24'b000000000000000000001000 : n28121_o;
  /* ../../HW/src/dp/dp_gen.vhd:1410:35  */
  assign n28125_o = src_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1411:41  */
  assign n28126_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1411:44  */
  assign n28128_o = n28126_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1413:44  */
  assign n28129_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1413:47  */
  assign n28131_o = n28129_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1413:22  */
  assign n28134_o = n28131_o ? 24'b000000000000000000100000 : 24'b000000000000010000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1411:22  */
  assign n28136_o = n28128_o ? 24'b000000000000000000000100 : n28134_o;
  /* ../../HW/src/dp/dp_gen.vhd:1418:35  */
  assign n28138_o = src_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1419:41  */
  assign n28139_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1419:44  */
  assign n28141_o = n28139_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1421:44  */
  assign n28142_o = src_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1421:47  */
  assign n28144_o = n28142_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1421:22  */
  assign n28147_o = n28144_o ? 24'b000000000000000000010000 : 24'b000000000000001000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1419:22  */
  assign n28149_o = n28141_o ? 24'b000000000000000000000010 : n28147_o;
  /* ../../HW/src/dp/dp_gen.vhd:1427:62  */
  assign n28150_o = n26310_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1418:19  */
  assign n28151_o = n28138_o ? n28149_o : n28150_o;
  /* ../../HW/src/dp/dp_gen.vhd:1410:19  */
  assign n28152_o = n28125_o ? n28136_o : n28151_o;
  /* ../../HW/src/dp/dp_gen.vhd:1402:19  */
  assign n28153_o = n28112_o ? n28123_o : n28152_o;
  /* ../../HW/src/dp/dp_gen.vhd:1431:60  */
  assign n28155_o = n28153_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1430:19  */
  assign n28156_o = source_double_precision ? n28155_o : n28153_o;
  /* ../../HW/src/dp/dp_gen.vhd:1436:63  */
  assign n28157_o = n26311_o[23:0];
  /* ../../HW/src/dp/dp_gen.vhd:1437:69  */
  assign n28158_o = n26311_o[47:24];
  /* ../../HW/src/dp/dp_gen.vhd:1438:67  */
  assign n28159_o = n26311_o[72:48];
  /* ../../HW/src/dp/dp_gen.vhd:1439:63  */
  assign n28160_o = n26311_o[121:98];
  /* ../../HW/src/dp/dp_gen.vhd:1440:69  */
  assign n28161_o = n26311_o[145:122];
  /* ../../HW/src/dp/dp_gen.vhd:1441:67  */
  assign n28162_o = n26311_o[170:146];
  /* ../../HW/src/dp/dp_gen.vhd:1442:63  */
  assign n28163_o = n26311_o[219:196];
  /* ../../HW/src/dp/dp_gen.vhd:1443:69  */
  assign n28164_o = n26311_o[243:220];
  /* ../../HW/src/dp/dp_gen.vhd:1444:67  */
  assign n28165_o = n26311_o[268:244];
  /* ../../HW/src/dp/dp_gen.vhd:1445:63  */
  assign n28166_o = n26311_o[317:294];
  /* ../../HW/src/dp/dp_gen.vhd:1446:69  */
  assign n28167_o = n26311_o[341:318];
  /* ../../HW/src/dp/dp_gen.vhd:1447:67  */
  assign n28168_o = n26311_o[366:342];
  /* ../../HW/src/dp/dp_gen.vhd:1448:63  */
  assign n28169_o = n26311_o[415:392];
  /* ../../HW/src/dp/dp_gen.vhd:1449:69  */
  assign n28170_o = n26311_o[439:416];
  /* ../../HW/src/dp/dp_gen.vhd:1450:67  */
  assign n28171_o = n26311_o[464:440];
  /* ../../HW/src/dp/dp_gen.vhd:1451:59  */
  assign n28172_o = n26311_o[624:593];
  /* ../../HW/src/dp/dp_gen.vhd:1452:63  */
  assign n28173_o = n26311_o[751:728];
  /* ../../HW/src/dp/dp_gen.vhd:1454:56  */
  assign n28174_o = n26311_o[564:540];
  /* ../../HW/src/dp/dp_gen.vhd:1455:65  */
  assign n28175_o = n26311_o[564:540];
  /* ../../HW/src/dp/dp_gen.vhd:1456:66  */
  assign n28176_o = n26311_o[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1457:71  */
  assign n28177_o = n26311_o[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1458:69  */
  assign n28178_o = n26311_o[775:752];
  /* ../../HW/src/dp/dp_gen.vhd:1460:32  */
  assign n28180_o = dst_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1461:126  */
  assign n28181_o = n26311_o[648:628];
  /* ../../HW/src/dp/dp_gen.vhd:1463:35  */
  assign n28184_o = dst_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1464:128  */
  assign n28185_o = n26311_o[648:627];
  /* ../../HW/src/dp/dp_gen.vhd:1466:35  */
  assign n28188_o = dst_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1467:128  */
  assign n28189_o = n26311_o[648:626];
  /* ../../HW/src/dp/dp_gen.vhd:1470:64  */
  assign n28191_o = n26311_o[648:625];
  assign n28192_o = {1'b0, n28189_o};
  /* ../../HW/src/dp/dp_gen.vhd:1466:19  */
  assign n28193_o = n28188_o ? n28192_o : n28191_o;
  assign n28194_o = {2'b00, n28185_o};
  /* ../../HW/src/dp/dp_gen.vhd:1463:19  */
  assign n28195_o = n28184_o ? n28194_o : n28193_o;
  assign n28196_o = {3'b000, n28181_o};
  /* ../../HW/src/dp/dp_gen.vhd:1460:19  */
  assign n28197_o = n28180_o ? n28196_o : n28195_o;
  /* ../../HW/src/dp/dp_gen.vhd:1473:42  */
  assign n28198_o = n26311_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1473:53  */
  assign n28200_o = n28198_o == 24'b000000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1473:19  */
  assign n28203_o = n28200_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1479:32  */
  assign n28205_o = dst_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1480:41  */
  assign n28206_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1480:44  */
  assign n28208_o = n28206_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1482:44  */
  assign n28210_o = dst_is_scatter_r[1:0];
  /* ../../HW/src/dp/dp_gen.vhd:1482:47  */
  assign n28212_o = n28210_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1482:22  */
  assign n28215_o = n28212_o ? 24'b000000000000000001000000 : 24'b000000000000100000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1480:22  */
  assign n28216_o = n28208_o ? 24'b000000000000000000001000 : n28215_o;
  /* ../../HW/src/dp/dp_gen.vhd:1487:35  */
  assign n28218_o = dst_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1488:41  */
  assign n28219_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1488:44  */
  assign n28221_o = n28219_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1490:44  */
  assign n28223_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1490:47  */
  assign n28225_o = n28223_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1490:22  */
  assign n28228_o = n28225_o ? 24'b000000000000000000100000 : 24'b000000000000010000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1488:22  */
  assign n28229_o = n28221_o ? 24'b000000000000000000000100 : n28228_o;
  /* ../../HW/src/dp/dp_gen.vhd:1495:35  */
  assign n28231_o = dst_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1496:41  */
  assign n28232_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1496:44  */
  assign n28234_o = n28232_o == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1498:44  */
  assign n28236_o = dst_is_scatter_r[3:2];
  /* ../../HW/src/dp/dp_gen.vhd:1498:47  */
  assign n28238_o = n28236_o == 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1498:22  */
  assign n28241_o = n28238_o ? 24'b000000000000000000010000 : 24'b000000000000001000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1496:22  */
  assign n28242_o = n28234_o ? 24'b000000000000000000000010 : n28241_o;
  /* ../../HW/src/dp/dp_gen.vhd:1504:70  */
  assign n28243_o = n26311_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1495:19  */
  assign n28244_o = n28231_o ? n28242_o : n28243_o;
  /* ../../HW/src/dp/dp_gen.vhd:1487:19  */
  assign n28245_o = n28218_o ? n28229_o : n28244_o;
  /* ../../HW/src/dp/dp_gen.vhd:1479:19  */
  assign n28246_o = n28205_o ? n28216_o : n28245_o;
  /* ../../HW/src/dp/dp_gen.vhd:1515:48  */
  assign n28248_o = instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1515:19  */
  assign n28250_o = n28248_o ? 1'b0 : instruction_stream_process_in;
  /* ../../HW/src/dp/dp_gen.vhd:1515:19  */
  assign n28252_o = n28248_o ? instruction_stream_process_in : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1526:50  */
  assign n28254_o = instruction_bus_id_source_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1526:102  */
  assign n28256_o = instruction_bus_id_dest_in == 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1526:72  */
  assign n28257_o = n28256_o & n28254_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:47  */
  assign n28258_o = n26310_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:1527:63  */
  assign n28259_o = ~n28258_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:92  */
  assign n28260_o = n26311_o[673];
  /* ../../HW/src/dp/dp_gen.vhd:1527:108  */
  assign n28261_o = ~n28260_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:68  */
  assign n28262_o = n28261_o & n28259_o;
  /* ../../HW/src/dp/dp_gen.vhd:1527:22  */
  assign n28265_o = n28262_o ? 2'b00 : 2'b01;
  /* ../../HW/src/dp/dp_gen.vhd:1532:78  */
  assign n28266_o = ~dest_double_precision;
  /* ../../HW/src/dp/dp_gen.vhd:1532:53  */
  assign n28267_o = n28266_o & source_double_precision;
  /* ../../HW/src/dp/dp_gen.vhd:1534:48  */
  assign n28268_o = ~source_double_precision;
  /* ../../HW/src/dp/dp_gen.vhd:1534:53  */
  assign n28269_o = dest_double_precision & n28268_o;
  /* ../../HW/src/dp/dp_gen.vhd:1534:19  */
  assign n28272_o = n28269_o ? 2'b10 : 2'b00;
  /* ../../HW/src/dp/dp_gen.vhd:1532:19  */
  assign n28274_o = n28267_o ? 2'b01 : n28272_o;
  /* ../../HW/src/dp/dp_gen.vhd:1526:19  */
  assign n28275_o = n28257_o ? n28265_o : n28274_o;
  /* ../../HW/src/dp/dp_gen.vhd:1543:32  */
  assign n28277_o = dst_vector == 3'b111;
  /* ../../HW/src/dp/dp_gen.vhd:1545:105  */
  assign n28279_o = instruction_gen_len_in[23:3];
  /* ../../HW/src/dp/dp_gen.vhd:1545:150  */
  assign n28281_o = n28279_o - 21'b000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1546:35  */
  assign n28283_o = dst_vector == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1548:107  */
  assign n28285_o = instruction_gen_len_in[23:2];
  /* ../../HW/src/dp/dp_gen.vhd:1548:154  */
  assign n28287_o = n28285_o - 22'b0000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1549:35  */
  assign n28289_o = dst_vector == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1551:107  */
  assign n28291_o = instruction_gen_len_in[23:1];
  /* ../../HW/src/dp/dp_gen.vhd:1551:154  */
  assign n28293_o = n28291_o - 23'b00000000000000000000001;
  /* ../../HW/src/dp/dp_gen.vhd:1553:58  */
  assign n28295_o = instruction_gen_len_in - 24'b000000000000000000000001;
  assign n28296_o = {1'b0, n28293_o};
  /* ../../HW/src/dp/dp_gen.vhd:1549:19  */
  assign n28297_o = n28289_o ? n28296_o : n28295_o;
  assign n28298_o = {2'b00, n28287_o};
  /* ../../HW/src/dp/dp_gen.vhd:1546:19  */
  assign n28299_o = n28283_o ? n28298_o : n28297_o;
  assign n28300_o = {3'b000, n28281_o};
  /* ../../HW/src/dp/dp_gen.vhd:1543:19  */
  assign n28301_o = n28277_o ? n28300_o : n28299_o;
  /* ../../HW/src/dp/dp_gen.vhd:1557:42  */
  assign n28303_o = n28301_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1557:19  */
  assign n28306_o = n28303_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1572:52  */
  assign n28307_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1573:52  */
  assign n28308_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1572:91  */
  assign n28309_o = {n28307_o, n28308_o};
  /* ../../HW/src/dp/dp_gen.vhd:1574:52  */
  assign n28310_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1573:80  */
  assign n28311_o = {n28309_o, n28310_o};
  /* ../../HW/src/dp/dp_gen.vhd:1575:52  */
  assign n28312_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1574:91  */
  assign n28313_o = {n28311_o, n28312_o};
  /* ../../HW/src/dp/dp_gen.vhd:1576:52  */
  assign n28314_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1575:80  */
  assign n28315_o = {n28313_o, n28314_o};
  /* ../../HW/src/dp/dp_gen.vhd:1577:52  */
  assign n28316_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1576:91  */
  assign n28317_o = {n28315_o, n28316_o};
  /* ../../HW/src/dp/dp_gen.vhd:1578:52  */
  assign n28318_o = instruction_data_in[15:8];
  /* ../../HW/src/dp/dp_gen.vhd:1577:80  */
  assign n28319_o = {n28317_o, n28318_o};
  /* ../../HW/src/dp/dp_gen.vhd:1579:52  */
  assign n28320_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1578:91  */
  assign n28321_o = {n28319_o, n28320_o};
  /* ../../HW/src/dp/dp_gen.vhd:1581:52  */
  assign n28322_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1582:52  */
  assign n28323_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1581:78  */
  assign n28324_o = {n28322_o, n28323_o};
  /* ../../HW/src/dp/dp_gen.vhd:1583:52  */
  assign n28325_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1582:78  */
  assign n28326_o = {n28324_o, n28325_o};
  /* ../../HW/src/dp/dp_gen.vhd:1584:52  */
  assign n28327_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1583:78  */
  assign n28328_o = {n28326_o, n28327_o};
  /* ../../HW/src/dp/dp_gen.vhd:1585:52  */
  assign n28329_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1584:78  */
  assign n28330_o = {n28328_o, n28329_o};
  /* ../../HW/src/dp/dp_gen.vhd:1586:52  */
  assign n28331_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1585:78  */
  assign n28332_o = {n28330_o, n28331_o};
  /* ../../HW/src/dp/dp_gen.vhd:1587:52  */
  assign n28333_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1586:78  */
  assign n28334_o = {n28332_o, n28333_o};
  /* ../../HW/src/dp/dp_gen.vhd:1588:52  */
  assign n28335_o = instruction_data_in[7:0];
  /* ../../HW/src/dp/dp_gen.vhd:1587:78  */
  assign n28336_o = {n28334_o, n28335_o};
  /* ../../HW/src/dp/dp_gen.vhd:1571:19  */
  assign n28337_o = source_double_precision ? n28321_o : n28336_o;
  /* ../../HW/src/dp/dp_gen.vhd:1592:44  */
  assign n28338_o = n26310_o[672:649];
  /* ../../HW/src/dp/dp_gen.vhd:1592:55  */
  assign n28340_o = n28338_o == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1592:19  */
  assign n28343_o = n28340_o ? 1'b1 : 1'b0;
  assign n28344_o = {n28067_o, n28076_o, n28073_o, n28070_o, n28066_o, n28065_o, n28064_o, n28063_o, n28062_o, n28061_o, n28060_o, n28059_o, n28058_o, n28057_o, n28056_o, n28055_o, n28054_o, n28053_o, n28052_o, n28051_o, n28050_o, n28049_o, n28048_o, n28047_o};
  assign n28345_o = {n28153_o, n28099_o, n28079_o, n28104_o};
  assign n28346_o = {n28080_o, n28078_o};
  assign n28354_o = {n28159_o, n28158_o, n28157_o};
  assign n28355_o = {n28162_o, n28161_o, n28160_o};
  assign n28356_o = {n28165_o, n28164_o, n28163_o};
  assign n28357_o = {n28168_o, n28167_o, n28166_o};
  assign n28358_o = {n28171_o, n28170_o, n28169_o};
  assign n28359_o = {n28176_o, n28175_o};
  assign n28360_o = {n28246_o, n28197_o, n28172_o};
  assign n28361_o = {n28178_o, n28173_o};
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n28380_o = instruction_latch_in ? n28174_o : d_burst_max_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n28381_o = instruction_latch_in ? n28301_o : currlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n28392_o = instruction_latch_in ? n28343_o : eof_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n28393_o = instruction_latch_in ? n28306_o : done_r;
  /* ../../HW/src/dp/dp_gen.vhd:1346:16  */
  assign n28411_o = instruction_latch_in ? n28104_o : n28032_burst_min_v;
  /* ../../HW/src/dp/dp_gen.vhd:1614:54  */
  assign n28414_o = n26310_o[97:73];
  /* ../../HW/src/dp/dp_gen.vhd:1615:54  */
  assign n28415_o = n26310_o[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1616:54  */
  assign n28416_o = n26310_o[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1617:54  */
  assign n28417_o = n26310_o[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1618:54  */
  assign n28418_o = n26310_o[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1638:40  */
  assign n28420_o = currlen_new == 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1638:16  */
  assign n28423_o = n28420_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1643:34  */
  assign n28424_o = ~s_burstlen_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1647:31  */
  assign n28425_o = ~s_i4_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1652:63  */
  assign n28426_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1654:31  */
  assign n28427_o = ~s_i3_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1661:63  */
  assign n28428_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1662:59  */
  assign n28429_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1664:31  */
  assign n28430_o = ~s_i2_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1673:63  */
  assign n28431_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1674:59  */
  assign n28432_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1675:59  */
  assign n28433_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1677:31  */
  assign n28434_o = ~s_i1_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1689:63  */
  assign n28435_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1690:59  */
  assign n28436_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1691:59  */
  assign n28437_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1692:59  */
  assign n28438_o = s_template_r[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1694:31  */
  assign n28439_o = ~s_i0_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1708:63  */
  assign n28440_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1709:59  */
  assign n28441_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1710:59  */
  assign n28442_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1711:59  */
  assign n28443_o = s_template_r[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1712:59  */
  assign n28444_o = s_template_r[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1715:28  */
  assign n28445_o = ~repeat_r;
  /* ../../HW/src/dp/dp_gen.vhd:1728:63  */
  assign n28446_o = s_template_r[592:568];
  /* ../../HW/src/dp/dp_gen.vhd:1729:59  */
  assign n28447_o = s_template_r[489:465];
  /* ../../HW/src/dp/dp_gen.vhd:1730:59  */
  assign n28448_o = s_template_r[391:367];
  /* ../../HW/src/dp/dp_gen.vhd:1731:59  */
  assign n28449_o = s_template_r[293:269];
  /* ../../HW/src/dp/dp_gen.vhd:1732:59  */
  assign n28450_o = s_template_r[195:171];
  /* ../../HW/src/dp/dp_gen.vhd:1733:59  */
  assign n28451_o = s_template_r[97:73];
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28453_o = n28439_o ? s_i0_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28455_o = n28439_o ? s_i0_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28456_o = n28439_o ? s_i0_start_new : n28451_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28457_o = n28439_o ? n28444_o : n28450_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28458_o = n28439_o ? n28443_o : n28449_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28459_o = n28439_o ? n28442_o : n28448_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28460_o = n28439_o ? n28441_o : n28447_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28461_o = n28439_o ? n28440_o : n28446_o;
  /* ../../HW/src/dp/dp_gen.vhd:1694:16  */
  assign n28462_o = n28439_o ? eof_r : n28445_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28463_o = n28434_o ? s_i0_r : n28453_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28465_o = n28434_o ? s_i1_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28466_o = n28434_o ? s_i0_count_r : n28455_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28468_o = n28434_o ? s_i1_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28469_o = n28434_o ? s_i0_start_r : n28456_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28470_o = n28434_o ? s_i1_start_new : n28457_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28471_o = n28434_o ? n28438_o : n28458_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28472_o = n28434_o ? n28437_o : n28459_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28473_o = n28434_o ? n28436_o : n28460_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28474_o = n28434_o ? n28435_o : n28461_o;
  /* ../../HW/src/dp/dp_gen.vhd:1677:16  */
  assign n28475_o = n28434_o ? eof_r : n28462_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28476_o = n28430_o ? s_i0_r : n28463_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28477_o = n28430_o ? s_i1_r : n28465_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28479_o = n28430_o ? s_i2_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28480_o = n28430_o ? s_i0_count_r : n28466_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28481_o = n28430_o ? s_i1_count_r : n28468_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28483_o = n28430_o ? s_i2_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28484_o = n28430_o ? s_i0_start_r : n28469_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28485_o = n28430_o ? s_i1_start_r : n28470_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28486_o = n28430_o ? s_i2_start_new : n28471_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28487_o = n28430_o ? n28433_o : n28472_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28488_o = n28430_o ? n28432_o : n28473_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28489_o = n28430_o ? n28431_o : n28474_o;
  /* ../../HW/src/dp/dp_gen.vhd:1664:16  */
  assign n28490_o = n28430_o ? eof_r : n28475_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28491_o = n28427_o ? s_i0_r : n28476_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28492_o = n28427_o ? s_i1_r : n28477_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28493_o = n28427_o ? s_i2_r : n28479_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28495_o = n28427_o ? s_i3_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28496_o = n28427_o ? s_i0_count_r : n28480_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28497_o = n28427_o ? s_i1_count_r : n28481_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28498_o = n28427_o ? s_i2_count_r : n28483_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28500_o = n28427_o ? s_i3_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28501_o = n28427_o ? s_i0_start_r : n28484_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28502_o = n28427_o ? s_i1_start_r : n28485_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28503_o = n28427_o ? s_i2_start_r : n28486_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28504_o = n28427_o ? s_i3_start_new : n28487_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28505_o = n28427_o ? n28429_o : n28488_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28506_o = n28427_o ? n28428_o : n28489_o;
  /* ../../HW/src/dp/dp_gen.vhd:1654:16  */
  assign n28507_o = n28427_o ? eof_r : n28490_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28508_o = n28425_o ? s_i0_r : n28491_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28509_o = n28425_o ? s_i1_r : n28492_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28510_o = n28425_o ? s_i2_r : n28493_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28511_o = n28425_o ? s_i3_r : n28495_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28513_o = n28425_o ? s_i4_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28514_o = n28425_o ? s_i0_count_r : n28496_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28515_o = n28425_o ? s_i1_count_r : n28497_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28516_o = n28425_o ? s_i2_count_r : n28498_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28517_o = n28425_o ? s_i3_count_r : n28500_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28519_o = n28425_o ? s_i4_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28520_o = n28425_o ? s_i0_start_r : n28501_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28521_o = n28425_o ? s_i1_start_r : n28502_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28522_o = n28425_o ? s_i2_start_r : n28503_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28523_o = n28425_o ? s_i3_start_r : n28504_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28524_o = n28425_o ? s_i4_start_new : n28505_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28525_o = n28425_o ? n28426_o : n28506_o;
  /* ../../HW/src/dp/dp_gen.vhd:1647:16  */
  assign n28526_o = n28425_o ? eof_r : n28507_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28527_o = n28424_o ? s_i0_r : n28508_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28528_o = n28424_o ? s_i1_r : n28509_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28529_o = n28424_o ? s_i2_r : n28510_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28530_o = n28424_o ? s_i3_r : n28511_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28531_o = n28424_o ? s_i4_r : n28513_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28532_o = n28424_o ? s_i0_count_r : n28514_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28533_o = n28424_o ? s_i1_count_r : n28515_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28534_o = n28424_o ? s_i2_count_r : n28516_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28535_o = n28424_o ? s_i3_count_r : n28517_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28536_o = n28424_o ? s_i4_count_r : n28519_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28538_o = n28424_o ? s_burstlen_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28540_o = n28424_o ? s_burstpos_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28541_o = n28424_o ? s_i0_start_r : n28520_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28542_o = n28424_o ? s_i1_start_r : n28521_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28543_o = n28424_o ? s_i2_start_r : n28522_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28544_o = n28424_o ? s_i3_start_r : n28523_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28545_o = n28424_o ? s_i4_start_r : n28524_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28546_o = n28424_o ? s_burstpos_start_new : n28525_o;
  /* ../../HW/src/dp/dp_gen.vhd:1643:16  */
  assign n28547_o = n28424_o ? eof_r : n28526_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:34  */
  assign n28548_o = ~d_burstlen_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1738:31  */
  assign n28549_o = ~d_i4_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1743:36  */
  assign n28550_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1743:51  */
  assign n28552_o = n28550_o == 3'b100;
  /* ../../HW/src/dp/dp_gen.vhd:1744:59  */
  assign n28553_o = d_template_r[463:440];
  /* ../../HW/src/dp/dp_gen.vhd:1744:33  */
  assign n28554_o = $unsigned(d_i4_new2) > $unsigned(n28553_o);
  /* ../../HW/src/dp/dp_gen.vhd:1743:55  */
  assign n28555_o = n28554_o & n28552_o;
  /* ../../HW/src/dp/dp_gen.vhd:1745:53  */
  assign n28556_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1747:53  */
  assign n28557_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1743:19  */
  assign n28558_o = n28555_o ? n28556_o : n28557_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:31  */
  assign n28559_o = ~d_i3_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1757:36  */
  assign n28561_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1757:51  */
  assign n28563_o = n28561_o == 3'b011;
  /* ../../HW/src/dp/dp_gen.vhd:1758:59  */
  assign n28564_o = d_template_r[365:342];
  /* ../../HW/src/dp/dp_gen.vhd:1758:33  */
  assign n28565_o = $unsigned(d_i3_new2) > $unsigned(n28564_o);
  /* ../../HW/src/dp/dp_gen.vhd:1757:55  */
  assign n28566_o = n28565_o & n28563_o;
  /* ../../HW/src/dp/dp_gen.vhd:1759:53  */
  assign n28567_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1761:53  */
  assign n28568_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1757:19  */
  assign n28569_o = n28566_o ? n28567_o : n28568_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:31  */
  assign n28570_o = ~d_i2_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1773:36  */
  assign n28572_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1773:51  */
  assign n28574_o = n28572_o == 3'b010;
  /* ../../HW/src/dp/dp_gen.vhd:1774:59  */
  assign n28575_o = d_template_r[267:244];
  /* ../../HW/src/dp/dp_gen.vhd:1774:33  */
  assign n28576_o = $unsigned(d_i2_new2) > $unsigned(n28575_o);
  /* ../../HW/src/dp/dp_gen.vhd:1773:55  */
  assign n28577_o = n28576_o & n28574_o;
  /* ../../HW/src/dp/dp_gen.vhd:1775:53  */
  assign n28578_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1777:53  */
  assign n28579_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1773:19  */
  assign n28580_o = n28577_o ? n28578_o : n28579_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:31  */
  assign n28581_o = ~d_i1_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1791:36  */
  assign n28583_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1791:51  */
  assign n28585_o = n28583_o == 3'b001;
  /* ../../HW/src/dp/dp_gen.vhd:1792:59  */
  assign n28586_o = d_template_r[169:146];
  /* ../../HW/src/dp/dp_gen.vhd:1792:33  */
  assign n28587_o = $unsigned(d_i1_new2) > $unsigned(n28586_o);
  /* ../../HW/src/dp/dp_gen.vhd:1791:55  */
  assign n28588_o = n28587_o & n28585_o;
  /* ../../HW/src/dp/dp_gen.vhd:1793:52  */
  assign n28589_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1795:52  */
  assign n28590_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1791:19  */
  assign n28591_o = n28588_o ? n28589_o : n28590_o;
  /* ../../HW/src/dp/dp_gen.vhd:1797:31  */
  assign n28592_o = ~d_i0_wrap;
  /* ../../HW/src/dp/dp_gen.vhd:1811:36  */
  assign n28594_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1811:51  */
  assign n28596_o = n28594_o == 3'b000;
  /* ../../HW/src/dp/dp_gen.vhd:1812:59  */
  assign n28597_o = d_template_r[71:48];
  /* ../../HW/src/dp/dp_gen.vhd:1812:33  */
  assign n28598_o = $unsigned(d_i0_new2) > $unsigned(n28597_o);
  /* ../../HW/src/dp/dp_gen.vhd:1811:55  */
  assign n28599_o = n28598_o & n28596_o;
  /* ../../HW/src/dp/dp_gen.vhd:1813:53  */
  assign n28600_o = d_template_r[539:515];
  /* ../../HW/src/dp/dp_gen.vhd:1815:53  */
  assign n28601_o = d_template_r[514:490];
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n28602_o = n28608_o ? n28600_o : n28601_o;
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n28605_o = n28592_o ? d_i0_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n28607_o = n28592_o ? d_i0_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1797:16  */
  assign n28608_o = n28599_o & n28592_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n28609_o = n28581_o ? d_i0_r : n28605_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n28611_o = n28581_o ? d_i1_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n28612_o = n28581_o ? d_i0_count_r : n28607_o;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n28614_o = n28581_o ? d_i1_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1779:16  */
  assign n28615_o = n28581_o ? n28591_o : n28602_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28616_o = n28570_o ? d_i0_r : n28609_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28617_o = n28570_o ? d_i1_r : n28611_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28619_o = n28570_o ? d_i2_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28620_o = n28570_o ? d_i0_count_r : n28612_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28621_o = n28570_o ? d_i1_count_r : n28614_o;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28623_o = n28570_o ? d_i2_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1763:16  */
  assign n28624_o = n28570_o ? n28580_o : n28615_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28625_o = n28559_o ? d_i0_r : n28616_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28626_o = n28559_o ? d_i1_r : n28617_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28627_o = n28559_o ? d_i2_r : n28619_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28629_o = n28559_o ? d_i3_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28630_o = n28559_o ? d_i0_count_r : n28620_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28631_o = n28559_o ? d_i1_count_r : n28621_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28632_o = n28559_o ? d_i2_count_r : n28623_o;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28634_o = n28559_o ? d_i3_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1749:16  */
  assign n28635_o = n28559_o ? n28569_o : n28624_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28636_o = n28549_o ? d_i0_r : n28625_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28637_o = n28549_o ? d_i1_r : n28626_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28638_o = n28549_o ? d_i2_r : n28627_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28639_o = n28549_o ? d_i3_r : n28629_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28641_o = n28549_o ? d_i4_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28642_o = n28549_o ? d_i0_count_r : n28630_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28643_o = n28549_o ? d_i1_count_r : n28631_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28644_o = n28549_o ? d_i2_count_r : n28632_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28645_o = n28549_o ? d_i3_count_r : n28634_o;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28647_o = n28549_o ? d_i4_count_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1738:16  */
  assign n28648_o = n28549_o ? n28558_o : n28635_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28649_o = n28548_o ? d_i0_r : n28636_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28650_o = n28548_o ? d_i1_r : n28637_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28651_o = n28548_o ? d_i2_r : n28638_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28652_o = n28548_o ? d_i3_r : n28639_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28653_o = n28548_o ? d_i4_r : n28641_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28654_o = n28548_o ? d_i0_count_r : n28642_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28655_o = n28548_o ? d_i1_count_r : n28643_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28656_o = n28548_o ? d_i2_count_r : n28644_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28657_o = n28548_o ? d_i3_count_r : n28645_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28658_o = n28548_o ? d_i4_count_r : n28647_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28659_o = n28548_o ? d_burst_max_r : n28648_o;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28661_o = n28548_o ? d_burstlen_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1735:16  */
  assign n28663_o = n28548_o ? d_burstpos_new : 24'b000000000000000000000000;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28665_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28667_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28669_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28671_o = reload ? 24'b000000000000000000000000 : n28527_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28673_o = reload ? 24'b000000000000000000000000 : n28528_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28675_o = reload ? 24'b000000000000000000000000 : n28529_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28677_o = reload ? 24'b000000000000000000000000 : n28530_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28679_o = reload ? 24'b000000000000000000000000 : n28531_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28681_o = reload ? 24'b000000000000000000000000 : n28532_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28683_o = reload ? 24'b000000000000000000000000 : n28533_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28685_o = reload ? 24'b000000000000000000000000 : n28534_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28687_o = reload ? 24'b000000000000000000000000 : n28535_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28689_o = reload ? 24'b000000000000000000000000 : n28536_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28691_o = reload ? 24'b000000000000000000000000 : n28538_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28693_o = reload ? 24'b000000000000000000000000 : n28540_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28694_o = reload ? n28414_o : n28541_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28695_o = reload ? n28415_o : n28542_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28696_o = reload ? n28416_o : n28543_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28697_o = reload ? n28417_o : n28544_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28698_o = reload ? n28418_o : n28545_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28699_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28700_o = reload ? n28411_o : n28546_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28702_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28704_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28706_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28708_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28710_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28712_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28714_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28716_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28718_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28720_o = reload ? 24'b000000000000000000000000 : n28649_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28722_o = reload ? 24'b000000000000000000000000 : n28650_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28724_o = reload ? 24'b000000000000000000000000 : n28651_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28726_o = reload ? 24'b000000000000000000000000 : n28652_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28728_o = reload ? 24'b000000000000000000000000 : n28653_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28730_o = reload ? 24'b000000000000000000000000 : n28654_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28732_o = reload ? 24'b000000000000000000000000 : n28655_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28734_o = reload ? 24'b000000000000000000000000 : n28656_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28736_o = reload ? 24'b000000000000000000000000 : n28657_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28738_o = reload ? 24'b000000000000000000000000 : n28658_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28739_o = reload ? n28380_o : n28659_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28741_o = reload ? 24'b000000000000000000000000 : n28661_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28743_o = reload ? 24'b000000000000000000000000 : n28663_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28744_o = reload ? n28381_o : currlen_new;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28747_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28748_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28749_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28750_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28751_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28752_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28753_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28754_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28755_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28756_o = reload ? n28392_o : n28547_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28757_o = reload ? n28393_o : n28423_o;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28758_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28759_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28760_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28761_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28762_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28763_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28764_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28765_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28766_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28767_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28768_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28769_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28770_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28771_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28772_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28773_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28774_o = instruction_latch_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28775_o = instruction_valid_in & reload;
  /* ../../HW/src/dp/dp_gen.vhd:1334:13  */
  assign n28777_o = reload ? n28046_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28782_o = n28665_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28784_o = n28667_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28786_o = n28669_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28804_o = n28699_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28807_o = n28702_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28809_o = n28704_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28811_o = n28706_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28813_o = n28708_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28815_o = n28710_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28817_o = n28712_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28819_o = n28714_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28821_o = n28716_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28823_o = n28718_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28839_o = reload & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28840_o = n28747_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28841_o = n28748_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28842_o = n28749_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28843_o = n28750_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28844_o = n28751_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28845_o = n28752_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28846_o = n28753_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28847_o = n28754_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28848_o = n28755_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28851_o = n28758_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28852_o = n28759_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28853_o = n28760_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28854_o = n28761_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28855_o = n28762_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28856_o = n28763_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28857_o = n28764_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28858_o = n28765_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28859_o = n28766_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28860_o = n28767_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28861_o = n28768_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28862_o = n28769_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28863_o = n28770_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28864_o = n28771_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28865_o = n28772_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28866_o = n28773_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28867_o = n28774_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28868_o = n28775_o & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28870_o = n28042_o ? n28777_o : 1'b0;
  /* ../../HW/src/dp/dp_gen.vhd:1333:10  */
  assign n28872_o = reload & n28042_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29125_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29126_o = n28872_o & n29125_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29127_o = n29126_o ? n28411_o : n28032_burst_min_v;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29128_q <= n29127_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29137_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29138_o = n28786_o & n29137_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29139_o = s_template_r[775:728];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29140_o = n29138_o ? n28346_o : n29139_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29141_q <= n29140_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29142_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29143_o = n28784_o & n29142_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29144_o = s_template_r[672:568];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29145_o = n29143_o ? n28345_o : n29144_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29146_q <= n29145_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29147_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29148_o = n28782_o & n29147_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29149_o = s_template_r[514:0];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29150_o = n29148_o ? n28344_o : n29149_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29151_q <= n29150_o;
  assign n29154_o = {n29141_q, 55'bZ, n29146_q, 53'bZ, n29151_q};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29155_o = n28042_o ? n28671_o : s_i0_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29156_q <= 24'b000000000000000000000000;
    else
      n29156_q <= n29155_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29157_o = n28042_o ? n28673_o : s_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29158_q <= 24'b000000000000000000000000;
    else
      n29158_q <= n29157_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29159_o = n28042_o ? n28675_o : s_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29160_q <= 24'b000000000000000000000000;
    else
      n29160_q <= n29159_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29161_o = n28042_o ? n28677_o : s_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29162_q <= 24'b000000000000000000000000;
    else
      n29162_q <= n29161_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29163_o = n28042_o ? n28679_o : s_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29164_q <= 24'b000000000000000000000000;
    else
      n29164_q <= n29163_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29165_o = n28042_o ? n28681_o : s_i0_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29166_q <= 24'b000000000000000000000000;
    else
      n29166_q <= n29165_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29167_o = n28042_o ? n28683_o : s_i1_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29168_q <= 24'b000000000000000000000000;
    else
      n29168_q <= n29167_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29169_o = n28042_o ? n28685_o : s_i2_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29170_q <= 24'b000000000000000000000000;
    else
      n29170_q <= n29169_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29171_o = n28042_o ? n28687_o : s_i3_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29172_q <= 24'b000000000000000000000000;
    else
      n29172_q <= n29171_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29173_o = n28042_o ? n28689_o : s_i4_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29174_q <= 24'b000000000000000000000000;
    else
      n29174_q <= n29173_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29175_o = n28042_o ? n28691_o : s_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29176_q <= 24'b000000000000000000000000;
    else
      n29176_q <= n29175_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29177_o = n28042_o ? n28693_o : s_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29178_q <= 24'b000000000000000000000000;
    else
      n29178_q <= n29177_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29181_o = n27236_o ? n27334_o : s_burstremain_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29182_q <= 24'b111111111111111111111111;
    else
      n29182_q <= n29181_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29183_o = n27236_o ? n27345_o : s_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29184_q <= 1'b1;
    else
      n29184_q <= n29183_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29185_o = n28042_o ? n28694_o : s_i0_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29186_q <= 25'b0000000000000000000000000;
    else
      n29186_q <= n29185_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29187_o = n28042_o ? n28695_o : s_i1_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29188_q <= 25'b0000000000000000000000000;
    else
      n29188_q <= n29187_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29189_o = n28042_o ? n28696_o : s_i2_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29190_q <= 25'b0000000000000000000000000;
    else
      n29190_q <= n29189_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29191_o = n28042_o ? n28697_o : s_i3_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29192_q <= 25'b0000000000000000000000000;
    else
      n29192_q <= n29191_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29193_o = n28042_o ? n28698_o : s_i4_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29194_q <= 25'b0000000000000000000000000;
    else
      n29194_q <= n29193_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29195_o = n28804_o ? n28156_o : s_burstpos_stride_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29196_q <= 24'b000000000000000000000000;
    else
      n29196_q <= n29195_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29197_o = n28042_o ? n28700_o : s_burstpos_start_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29198_q <= 25'b0000000000000000000000000;
    else
      n29198_q <= n29197_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29199_o = n27236_o ? n27398_o : s_burstpos_start_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29200_q <= 4'b0000;
    else
      n29200_q <= n29199_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29201_o = n27236_o ? s_burstpos_start_rr : s_burstpos_start_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29202_q <= 4'b0000;
    else
      n29202_q <= n29201_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29203_o = n27236_o ? s_burstpos_start_rrr : s_burstpos_start_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29204_q <= 4'b0000;
    else
      n29204_q <= n29203_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29205_o = n27236_o ? n27287_o : s_burstpos_end_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29206_q <= 27'b000000000000000000000000000;
    else
      n29206_q <= n29205_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29207_o = n27236_o ? n27296_o : s_burstpos_end_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29208_q <= 4'b0000;
    else
      n29208_q <= n29207_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29209_o = n27236_o ? n27311_o : s_burstpos_end_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29210_q <= 4'b0000;
    else
      n29210_q <= n29209_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29211_o = n27236_o ? n27425_o : d_burstpos_end_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29212_q <= 27'b000000000000000000000000000;
    else
      n29212_q <= n29211_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29213_o = n27236_o ? n27434_o : d_burstpos_end_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29214_q <= 4'b0000;
    else
      n29214_q <= n29213_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29215_o = n27236_o ? n27449_o : d_burstpos_end_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29216_q <= 4'b0000;
    else
      n29216_q <= n29215_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29217_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29218_o = n28823_o & n29217_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29219_o = d_template_r[775:728];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29220_o = n29218_o ? n28361_o : n29219_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29221_q <= n29220_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29222_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29223_o = n28821_o & n29222_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29224_o = d_template_r[672:593];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29225_o = n29223_o ? n28360_o : n29224_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29226_q <= n29225_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29227_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29228_o = n28819_o & n29227_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29229_o = d_template_r[567:565];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29230_o = n29228_o ? n28177_o : n29229_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29231_q <= n29230_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29232_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29233_o = n28817_o & n29232_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29234_o = d_template_r[539:490];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29235_o = n29233_o ? n28359_o : n29234_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29236_q <= n29235_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29237_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29238_o = n28815_o & n29237_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29239_o = d_template_r[464:392];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29240_o = n29238_o ? n28358_o : n29239_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29241_q <= n29240_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29242_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29243_o = n28813_o & n29242_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29244_o = d_template_r[366:294];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29245_o = n29243_o ? n28357_o : n29244_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29246_q <= n29245_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29247_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29248_o = n28811_o & n29247_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29249_o = d_template_r[268:196];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29250_o = n29248_o ? n28356_o : n29249_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29251_q <= n29250_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29252_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29253_o = n28809_o & n29252_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29254_o = d_template_r[170:98];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29255_o = n29253_o ? n28355_o : n29254_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29256_q <= n29255_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29257_o = ~n28038_o;
  /* ../../HW/src/dp/dp_gen.vhd:1250:1  */
  assign n29258_o = n28807_o & n29257_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29259_o = d_template_r[72:0];
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29260_o = n29258_o ? n28354_o : n29259_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in)
    n29261_q <= n29260_o;
  assign n29270_o = {n29221_q, 55'bZ, n29226_q, 25'bZ, n29231_q, 25'bZ, n29236_q, 25'bZ, n29241_q, 25'bZ, n29246_q, 25'bZ, n29251_q, 25'bZ, n29256_q, 25'bZ, n29261_q};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29271_o = n28042_o ? n28720_o : d_i0_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29272_q <= 24'b000000000000000000000000;
    else
      n29272_q <= n29271_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29273_o = n28042_o ? n28722_o : d_i1_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29274_q <= 24'b000000000000000000000000;
    else
      n29274_q <= n29273_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29275_o = n28042_o ? n28724_o : d_i2_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29276_q <= 24'b000000000000000000000000;
    else
      n29276_q <= n29275_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29277_o = n28042_o ? n28726_o : d_i3_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29278_q <= 24'b000000000000000000000000;
    else
      n29278_q <= n29277_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29279_o = n28042_o ? n28728_o : d_i4_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29280_q <= 24'b000000000000000000000000;
    else
      n29280_q <= n29279_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29281_o = n28042_o ? n28730_o : d_i0_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29282_q <= 24'b000000000000000000000000;
    else
      n29282_q <= n29281_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29283_o = n28042_o ? n28732_o : d_i1_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29284_q <= 24'b000000000000000000000000;
    else
      n29284_q <= n29283_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29285_o = n28042_o ? n28734_o : d_i2_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29286_q <= 24'b000000000000000000000000;
    else
      n29286_q <= n29285_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29287_o = n28042_o ? n28736_o : d_i3_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29288_q <= 24'b000000000000000000000000;
    else
      n29288_q <= n29287_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29289_o = n28042_o ? n28738_o : d_i4_count_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29290_q <= 24'b000000000000000000000000;
    else
      n29290_q <= n29289_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29291_o = n28042_o ? n28739_o : d_burst_max_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29292_q <= 25'b0000000000000000000000000;
    else
      n29292_q <= n29291_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29293_o = n28042_o ? n28741_o : d_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29294_q <= 24'b000000000000000000000000;
    else
      n29294_q <= n29293_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29295_o = n28042_o ? n28743_o : d_burstpos_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29296_q <= 24'b000000000000000000000000;
    else
      n29296_q <= n29295_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29299_o = n27236_o ? n27472_o : d_burstremain_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29300_q <= 24'b111111111111111111111111;
    else
      n29300_q <= n29299_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29301_o = n27236_o ? n27477_o : d_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29302_q <= 1'b1;
    else
      n29302_q <= n29301_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29303_o = n28042_o ? n28744_o : currlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29304_q <= 24'b000000000000000000000000;
    else
      n29304_q <= n29303_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29307_o = n28839_o ? instruction_valid_in : running_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29308_q <= 1'b0;
    else
      n29308_q <= n29307_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29309_o = n27236_o ? running_r : running_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29310_q <= 1'b0;
    else
      n29310_q <= n29309_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29311_o = n27236_o ? running_rr : running_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29312_q <= 1'b0;
    else
      n29312_q <= n29311_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29313_o = n27236_o ? running_rrr : running_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29314_q <= 1'b0;
    else
      n29314_q <= n29313_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29315_o = n27236_o ? n27536_o : gen_valid_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29316_q <= 3'b000;
    else
      n29316_q <= n29315_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29317_o = n28840_o ? instruction_bus_id_dest_in : dp_dst_bus_id_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29318_q <= 2'b00;
    else
      n29318_q <= n29317_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29319_o = n27236_o ? dp_dst_bus_id_r : dp_dst_bus_id_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29320_q <= 2'b00;
    else
      n29320_q <= n29319_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29321_o = n27236_o ? dp_dst_bus_id_rr : dp_dst_bus_id_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29322_q <= 2'b00;
    else
      n29322_q <= n29321_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29323_o = n27236_o ? dp_dst_bus_id_rrr : dp_dst_bus_id_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29324_q <= 2'b00;
    else
      n29324_q <= n29323_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29325_o = n28841_o ? instruction_bus_id_source_in : dp_src_bus_id_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29326_q <= 2'b00;
    else
      n29326_q <= n29325_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29327_o = n27236_o ? dp_src_bus_id_r : dp_src_bus_id_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29328_q <= 2'b00;
    else
      n29328_q <= n29327_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29329_o = n27236_o ? dp_src_bus_id_rr : dp_src_bus_id_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29330_q <= 2'b00;
    else
      n29330_q <= n29329_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29331_o = n27236_o ? dp_src_bus_id_rrr : dp_src_bus_id_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29332_q <= 2'b00;
    else
      n29332_q <= n29331_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29333_o = n28842_o ? instruction_data_type_dest_in : dp_dst_data_type_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29334_q <= 2'b00;
    else
      n29334_q <= n29333_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29335_o = n27236_o ? dp_dst_data_type_r : dp_dst_data_type_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29336_q <= 2'b00;
    else
      n29336_q <= n29335_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29337_o = n27236_o ? dp_dst_data_type_rr : dp_dst_data_type_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29338_q <= 2'b00;
    else
      n29338_q <= n29337_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29339_o = n27236_o ? dp_dst_data_type_rrr : dp_dst_data_type_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29340_q <= 2'b00;
    else
      n29340_q <= n29339_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29341_o = n28843_o ? instruction_data_type_source_in : dp_src_data_type_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29342_q <= 2'b00;
    else
      n29342_q <= n29341_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29343_o = n27236_o ? dp_src_data_type_r : dp_src_data_type_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29344_q <= 2'b00;
    else
      n29344_q <= n29343_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29345_o = n27236_o ? dp_src_data_type_rr : dp_src_data_type_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29346_q <= 2'b00;
    else
      n29346_q <= n29345_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29347_o = n27236_o ? dp_src_data_type_rrr : dp_src_data_type_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29348_q <= 2'b00;
    else
      n29348_q <= n29347_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29349_o = n28844_o ? instruction_data_model_source_in : dp_src_data_model_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29350_q <= 2'b00;
    else
      n29350_q <= n29349_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29351_o = n27236_o ? dp_src_data_model_r : dp_src_data_model_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29352_q <= 2'b00;
    else
      n29352_q <= n29351_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29353_o = n27236_o ? dp_src_data_model_rr : dp_src_data_model_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29354_q <= 2'b00;
    else
      n29354_q <= n29353_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29355_o = n27236_o ? dp_src_data_model_rrr : dp_src_data_model_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29356_q <= 2'b00;
    else
      n29356_q <= n29355_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29357_o = n28845_o ? instruction_data_model_dest_in : dp_dst_data_model_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29358_q <= 2'b00;
    else
      n29358_q <= n29357_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29359_o = n27236_o ? dp_dst_data_model_r : dp_dst_data_model_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29360_q <= 2'b00;
    else
      n29360_q <= n29359_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29361_o = n27236_o ? dp_dst_data_model_rr : dp_dst_data_model_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29362_q <= 2'b00;
    else
      n29362_q <= n29361_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29363_o = n27236_o ? dp_dst_data_model_rrr : dp_dst_data_model_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29364_q <= 2'b00;
    else
      n29364_q <= n29363_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29365_o = n28846_o ? instruction_thread_in : dp_thread_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29366_q <= 1'b0;
    else
      n29366_q <= n29365_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29367_o = n27236_o ? dp_thread_r : dp_thread_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29368_q <= 1'b0;
    else
      n29368_q <= n29367_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29369_o = n27236_o ? dp_thread_rr : dp_thread_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29370_q <= 1'b0;
    else
      n29370_q <= n29369_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29371_o = n27236_o ? dp_thread_rrr : dp_thread_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29372_q <= 1'b0;
    else
      n29372_q <= n29371_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29373_o = n28847_o ? instruction_mcast_in : dp_mcast_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29374_q <= 6'b111111;
    else
      n29374_q <= n29373_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29375_o = n27236_o ? dp_mcast_r : dp_mcast_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29376_q <= 6'b111111;
    else
      n29376_q <= n29375_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29377_o = n27236_o ? dp_mcast_rr : dp_mcast_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29378_q <= 6'b111111;
    else
      n29378_q <= n29377_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29379_o = n27236_o ? dp_mcast_rrr : dp_mcast_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29380_q <= 6'b111111;
    else
      n29380_q <= n29379_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29381_o = n28848_o ? n28337_o : data_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29382_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n29382_q <= n29381_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29383_o = n27236_o ? data_r : data_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29384_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n29384_q <= n29383_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29385_o = n27236_o ? data_rr : data_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29386_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n29386_q <= n29385_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29387_o = n27236_o ? data_rrr : data_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29388_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n29388_q <= n29387_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29389_o = n27236_o ? n27254_o : s_bufsize_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29390_q <= 24'b000000000000000000000000;
    else
      n29390_q <= n29389_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29391_o = n27236_o ? s_bufsize_r : s_bufsize_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29392_q <= 24'b000000000000000000000000;
    else
      n29392_q <= n29391_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29393_o = n27236_o ? n27253_o : s_temp1_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29394_q <= 24'b000000000000000000000000;
    else
      n29394_q <= n29393_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29395_o = n27236_o ? n27255_o : s_temp2_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29396_q <= 32'b00000000000000000000000000000000;
    else
      n29396_q <= n29395_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29397_o = n27236_o ? n27257_o : s_temp3_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29398_q <= 24'b000000000000000000000000;
    else
      n29398_q <= n29397_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29399_o = n27236_o ? n27259_o : s_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29400_q <= 24'b000000000000000000000000;
    else
      n29400_q <= n29399_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29401_o = n27236_o ? n27260_o : s_temp5_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29402_q <= 24'b000000000000000000000000;
    else
      n29402_q <= n29401_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29403_o = n27236_o ? s_temp2_r : s_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29404_q <= 32'b00000000000000000000000000000000;
    else
      n29404_q <= n29403_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29405_o = n27236_o ? n27265_o : s_gen_addr_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29406_q <= 32'b00000000000000000000000000000000;
    else
      n29406_q <= n29405_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29407_o = n27236_o ? n27381_o : s_gen_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29408_q <= 5'b00000;
    else
      n29408_q <= n29407_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29409_o = n27236_o ? n27273_o : s_gen_burstlen_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29410_q <= 5'b00000;
    else
      n29410_q <= n29409_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29411_o = n27236_o ? n27278_o : s_gen_burstlen_progress_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29412_q <= 1'b0;
    else
      n29412_q <= n29411_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29413_o = n27236_o ? n27403_o : d_bufsize_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29414_q <= 24'b000000000000000000000000;
    else
      n29414_q <= n29413_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29415_o = n27236_o ? d_bufsize_r : d_bufsize_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29416_q <= 24'b000000000000000000000000;
    else
      n29416_q <= n29415_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29417_o = n27236_o ? n27405_o : d_temp1_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29418_q <= 24'b000000000000000000000000;
    else
      n29418_q <= n29417_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29419_o = n27236_o ? n27406_o : d_temp2_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29420_q <= 32'b00000000000000000000000000000000;
    else
      n29420_q <= n29419_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29421_o = n27236_o ? n27408_o : d_temp3_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29422_q <= 24'b000000000000000000000000;
    else
      n29422_q <= n29421_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29423_o = n27236_o ? n27410_o : d_temp4_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29424_q <= 24'b000000000000000000000000;
    else
      n29424_q <= n29423_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29425_o = n27236_o ? n27411_o : d_temp5_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29426_q <= 24'b000000000000000000000000;
    else
      n29426_q <= n29425_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29427_o = n27236_o ? d_temp2_r : d_temp4_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29428_q <= 32'b00000000000000000000000000000000;
    else
      n29428_q <= n29427_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29429_o = n27236_o ? n27416_o : d_gen_addr_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29430_q <= 32'b00000000000000000000000000000000;
    else
      n29430_q <= n29429_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29431_o = n27236_o ? n27513_o : d_gen_burstlen_r;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29432_q <= 5'b00000;
    else
      n29432_q <= n29431_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29433_o = n27236_o ? d_gen_burstlen_r : d_gen_burstlen_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29434_q <= 5'b00000;
    else
      n29434_q <= n29433_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29435_o = n28042_o ? n28756_o : eof_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29436_q <= 1'b0;
    else
      n29436_q <= n29435_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29437_o = n27236_o ? eof_r : eof_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29438_q <= 1'b0;
    else
      n29438_q <= n29437_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29439_o = n27236_o ? eof_rr : eof_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29440_q <= 1'b0;
    else
      n29440_q <= n29439_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29441_o = n27236_o ? eof_rrr : eof_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29442_q <= 1'b0;
    else
      n29442_q <= n29441_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29443_o = n28042_o ? n28757_o : done_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29444_q <= 1'b1;
    else
      n29444_q <= n29443_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29445_o = n28851_o ? instruction_repeat_in : repeat_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29446_q <= 1'b0;
    else
      n29446_q <= n29445_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29447_o = n28852_o ? n28275_o : data_flow_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29448_q <= 2'b00;
    else
      n29448_q <= n29447_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29449_o = n27236_o ? data_flow_r : data_flow_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29450_q <= 2'b00;
    else
      n29450_q <= n29449_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29451_o = n27236_o ? data_flow_rr : data_flow_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29452_q <= 2'b00;
    else
      n29452_q <= n29451_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29453_o = n27236_o ? data_flow_rrr : data_flow_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29454_q <= 2'b00;
    else
      n29454_q <= n29453_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29455_o = n28853_o ? n28250_o : stream_src_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29456_q <= 1'b0;
    else
      n29456_q <= n29455_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29457_o = n27236_o ? stream_src_r : stream_src_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29458_q <= 1'b0;
    else
      n29458_q <= n29457_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29459_o = n27236_o ? stream_src_rr : stream_src_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29460_q <= 1'b0;
    else
      n29460_q <= n29459_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29461_o = n27236_o ? stream_src_rrr : stream_src_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29462_q <= 1'b0;
    else
      n29462_q <= n29461_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29463_o = n28854_o ? n28252_o : stream_dest_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29464_q <= 1'b0;
    else
      n29464_q <= n29463_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29465_o = n27236_o ? stream_dest_r : stream_dest_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29466_q <= 1'b0;
    else
      n29466_q <= n29465_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29467_o = n27236_o ? stream_dest_rr : stream_dest_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29468_q <= 1'b0;
    else
      n29468_q <= n29467_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29469_o = n27236_o ? stream_dest_rrr : stream_dest_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29470_q <= 1'b0;
    else
      n29470_q <= n29469_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29471_o = n28855_o ? instruction_vm_in : vm_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29472_q <= 1'b0;
    else
      n29472_q <= n29471_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29473_o = n27236_o ? vm_r : vm_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29474_q <= 1'b0;
    else
      n29474_q <= n29473_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29475_o = n27236_o ? vm_rr : vm_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29476_q <= 1'b0;
    else
      n29476_q <= n29475_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29477_o = n27236_o ? vm_rrr : vm_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29478_q <= 1'b0;
    else
      n29478_q <= n29477_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29479_o = n28856_o ? instruction_stream_process_id_in : stream_id_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29480_q <= 2'b00;
    else
      n29480_q <= n29479_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29481_o = n27236_o ? stream_id_r : stream_id_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29482_q <= 2'b00;
    else
      n29482_q <= n29481_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29483_o = n27236_o ? stream_id_rr : stream_id_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29484_q <= 2'b00;
    else
      n29484_q <= n29483_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29485_o = n27236_o ? stream_id_rrr : stream_id_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29486_q <= 2'b00;
    else
      n29486_q <= n29485_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29487_o = n28857_o ? source_double_precision : src_double_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29488_q <= 1'b0;
    else
      n29488_q <= n29487_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29489_o = n27236_o ? src_double_r : src_double_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29490_q <= 1'b0;
    else
      n29490_q <= n29489_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29491_o = n27236_o ? src_double_rr : src_double_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29492_q <= 1'b0;
    else
      n29492_q <= n29491_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29495_o = n28858_o ? dest_double_precision : dst_double_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29496_q <= 1'b0;
    else
      n29496_q <= n29495_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29497_o = n27236_o ? dst_double_r : dst_double_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29498_q <= 1'b0;
    else
      n29498_q <= n29497_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29499_o = n27236_o ? dst_double_rr : dst_double_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29500_q <= 1'b0;
    else
      n29500_q <= n29499_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29503_o = n28859_o ? src_vector : src_vector_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29504_q <= 3'b000;
    else
      n29504_q <= n29503_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29505_o = n27236_o ? src_vector_r : src_vector_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29506_q <= 3'b000;
    else
      n29506_q <= n29505_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29507_o = n27236_o ? src_vector_rr : src_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29508_q <= 3'b000;
    else
      n29508_q <= n29507_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29509_o = n27236_o ? n27386_o : src_vector_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29510_q <= 3'b000;
    else
      n29510_q <= n29509_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29511_o = n28860_o ? dst_vector : dst_vector_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29512_q <= 3'b000;
    else
      n29512_q <= n29511_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29513_o = n27236_o ? dst_vector_r : dst_vector_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29514_q <= 3'b000;
    else
      n29514_q <= n29513_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29515_o = n27236_o ? dst_vector_rr : dst_vector_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29516_q <= 3'b000;
    else
      n29516_q <= n29515_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29517_o = n27236_o ? n27402_o : dst_vector_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29518_q <= 3'b000;
    else
      n29518_q <= n29517_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29519_o = n28861_o ? instruction_source_addr_mode_in : src_addr_mode_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29520_q <= 1'b0;
    else
      n29520_q <= n29519_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29521_o = n27236_o ? src_addr_mode_r : src_addr_mode_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29522_q <= 1'b0;
    else
      n29522_q <= n29521_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29523_o = n27236_o ? src_addr_mode_rr : src_addr_mode_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29524_q <= 1'b0;
    else
      n29524_q <= n29523_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29525_o = n27236_o ? src_addr_mode_rrr : src_addr_mode_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29526_q <= 1'b0;
    else
      n29526_q <= n29525_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29527_o = n28862_o ? instruction_dest_addr_mode_in : dst_addr_mode_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29528_q <= 1'b0;
    else
      n29528_q <= n29527_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29529_o = n27236_o ? dst_addr_mode_r : dst_addr_mode_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29530_q <= 1'b0;
    else
      n29530_q <= n29529_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29531_o = n27236_o ? dst_addr_mode_rr : dst_addr_mode_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29532_q <= 1'b0;
    else
      n29532_q <= n29531_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29533_o = n27236_o ? dst_addr_mode_rrr : dst_addr_mode_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29534_q <= 1'b0;
    else
      n29534_q <= n29533_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29535_o = n28863_o ? src_scatter : src_scatter_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29536_q <= 2'b00;
    else
      n29536_q <= n29535_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29537_o = n27236_o ? src_scatter_r : src_scatter_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29538_q <= 2'b00;
    else
      n29538_q <= n29537_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29539_o = n27236_o ? src_scatter_rr : src_scatter_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29540_q <= 2'b00;
    else
      n29540_q <= n29539_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29541_o = n27236_o ? src_scatter_rrr : src_scatter_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29542_q <= 2'b00;
    else
      n29542_q <= n29541_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29543_o = n28864_o ? dst_scatter : dst_scatter_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29544_q <= 2'b00;
    else
      n29544_q <= n29543_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29545_o = n27236_o ? dst_scatter_r : dst_scatter_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29546_q <= 2'b00;
    else
      n29546_q <= n29545_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29547_o = n27236_o ? dst_scatter_rr : dst_scatter_rrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29548_q <= 2'b00;
    else
      n29548_q <= n29547_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29549_o = n27236_o ? dst_scatter_rrr : dst_scatter_rrrr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29550_q <= 2'b00;
    else
      n29550_q <= n29549_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29551_o = n28865_o ? n28110_o : src_is_burst_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29552_q <= 1'b0;
    else
      n29552_q <= n29551_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29553_o = n27236_o ? src_is_burst_r : src_is_burst_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29554_q <= 1'b0;
    else
      n29554_q <= n29553_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29555_o = n28866_o ? n28203_o : dst_is_burst_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29556_q <= 1'b0;
    else
      n29556_q <= n29555_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  assign n29557_o = n27236_o ? dst_is_burst_r : dst_is_burst_rr;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29558_q <= 1'b0;
    else
      n29558_q <= n29557_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n26394_o)
    if (n26394_o)
      n29560_q <= 3'b000;
    else
      n29560_q <= n26855_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n26394_o)
    if (n26394_o)
      n29561_q <= 3'b000;
    else
      n29561_q <= n26857_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n26394_o)
    if (n26394_o)
      n29562_q <= 6'b000000;
    else
      n29562_q <= n26859_o;
  /* ../../HW/src/dp/dp_gen.vhd:537:1  */
  always @(posedge clock_in or posedge n26394_o)
    if (n26394_o)
      n29563_q <= 6'b000000;
    else
      n29563_q <= n26861_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29564_o = n28867_o ? n28077_o : s_burst_actual_max_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29565_q <= 25'b0000000000000000000000000;
    else
      n29565_q <= n29564_o;
  /* ../../HW/src/dp/dp_gen.vhd:1256:4  */
  assign n29566_o = {14'b00000000000000, dest_double_precision, dst_scatter, dst_vector, instruction_bus_id_dest_in, source_double_precision, src_scatter, src_vector, instruction_bus_id_source_in, 2'b01};
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  assign n29567_o = n28868_o ? log : log_r;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29568_q <= 32'b00000000000000000000000000000000;
    else
      n29568_q <= n29567_o;
  /* ../../HW/src/dp/dp_gen.vhd:1331:7  */
  always @(posedge clock_in or posedge n28038_o)
    if (n28038_o)
      n29569_q <= 1'b0;
    else
      n29569_q <= n28870_o;
  /* ../../HW/src/dp/dp_gen.vhd:914:9  */
  always @(posedge clock_in or posedge n27234_o)
    if (n27234_o)
      n29572_q <= 1'b0;
    else
      n29572_q <= n27632_o;
  /* ../../HW/src/dp/dp_gen.vhd:121:16  */
  assign n29573_o = wr_full_in[0];
  /* ../../HW/src/dp/dp_gen.vhd:120:16  */
  assign n29574_o = wr_full_in[1];
  /* ../../HW/src/dp/dp_gen.vhd:116:16  */
  assign n29575_o = wr_full_in[2];
  /* ../../HW/src/dp/dp_gen.vhd:115:16  */
  assign n29576_o = dp_dst_bus_id_rrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:926:46  */
  assign n29577_o = n29576_o ? n29574_o : n29573_o;
  /* ../../HW/src/dp/dp_gen.vhd:113:16  */
  assign n29578_o = dp_dst_bus_id_rrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:926:46  */
  assign n29579_o = n29578_o ? n29575_o : n29577_o;
  /* ../../HW/src/dp/dp_gen.vhd:926:46  */
  assign n29580_o = wr_maxburstlen_in[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:926:47  */
  assign n29581_o = wr_maxburstlen_in[9:5];
  /* ../../HW/src/dp/dp_gen.vhd:111:16  */
  assign n29582_o = wr_maxburstlen_in[14:10];
  /* ../../HW/src/dp/dp_gen.vhd:110:16  */
  assign n29583_o = dp_dst_bus_id_rrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:985:56  */
  assign n29584_o = n29583_o ? n29581_o : n29580_o;
  /* ../../HW/src/dp/dp_gen.vhd:108:16  */
  assign n29585_o = dp_dst_bus_id_rrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:985:56  */
  assign n29586_o = n29585_o ? n29582_o : n29584_o;
  /* ../../HW/src/dp/dp_gen.vhd:985:56  */
  assign n29587_o = wr_maxburstlen_in[4:0];
  /* ../../HW/src/dp/dp_gen.vhd:985:57  */
  assign n29588_o = wr_maxburstlen_in[9:5];
  /* ../../HW/src/dp/dp_gen.vhd:106:16  */
  assign n29589_o = wr_maxburstlen_in[14:10];
  /* ../../HW/src/dp/dp_gen.vhd:105:16  */
  assign n29590_o = dp_dst_bus_id_rrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:986:54  */
  assign n29591_o = n29590_o ? n29588_o : n29587_o;
  /* ../../HW/src/dp/dp_gen.vhd:103:16  */
  assign n29592_o = dp_dst_bus_id_rrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:986:54  */
  assign n29593_o = n29592_o ? n29589_o : n29591_o;
  /* ../../HW/src/dp/dp_gen.vhd:986:54  */
  assign n29594_o = wr_full_in[0];
  /* ../../HW/src/dp/dp_gen.vhd:986:55  */
  assign n29595_o = wr_full_in[1];
  /* ../../HW/src/dp/dp_gen.vhd:101:16  */
  assign n29596_o = wr_full_in[2];
  /* ../../HW/src/dp/dp_gen.vhd:100:16  */
  assign n29597_o = dp_dst_bus_id_rrrr[0];
  /* ../../HW/src/dp/dp_gen.vhd:1240:46  */
  assign n29598_o = n29597_o ? n29595_o : n29594_o;
  /* ../../HW/src/dp/dp_gen.vhd:98:16  */
  assign n29599_o = dp_dst_bus_id_rrrr[1];
  /* ../../HW/src/dp/dp_gen.vhd:1240:46  */
  assign n29600_o = n29599_o ? n29596_o : n29598_o;
endmodule

module scfifo_67_8_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [66:0] data_in,
   input  write_in,
   input  read_in,
   output [66:0] q_out,
   output [7:0] ravail_out,
   output [7:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [66:0] q;
  wire [7:0] address_a;
  wire [7:0] address_b;
  wire [7:0] waddr_r;
  wire [7:0] waddr_rr;
  wire [7:0] raddr_r;
  wire [7:0] raddr;
  wire [7:0] ravail;
  wire [7:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [66:0] ram_i_n26242;
  wire [66:0] ram_i_q_b;
  wire [7:0] n26245_o;
  wire [7:0] n26246_o;
  wire n26247_o;
  wire n26250_o;
  wire n26251_o;
  wire [7:0] n26254_o;
  wire [7:0] n26255_o;
  wire n26258_o;
  wire [7:0] n26261_o;
  wire [7:0] n26263_o;
  wire n26264_o;
  wire n26267_o;
  wire [7:0] n26269_o;
  wire n26270_o;
  wire n26273_o;
  wire n26275_o;
  wire n26277_o;
  wire n26280_o;
  wire [7:0] n26302_o;
  reg [7:0] n26303_q;
  reg [7:0] n26304_q;
  reg [7:0] n26305_q;
  reg n26307_q;
  reg n26308_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n26247_o;
  assign full_out = full_r;
  assign almost_full_out = n26251_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n26242; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n26303_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n26304_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n26305_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n26255_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n26245_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n26246_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n26307_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n26308_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n26242 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_256_256_8_8_67_67 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n26245_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n26246_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n26247_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n26250_o = $unsigned(wused) >= $unsigned(8'b00000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n26251_o = n26250_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n26254_o = raddr_r + 8'b00000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n26255_o = read_in ? n26254_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n26258_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n26261_o = waddr_r + 8'b00000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n26263_o = waddr_r + 8'b00000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n26264_o = n26263_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n26267_o = n26264_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n26269_o = waddr_r + 8'b00000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n26270_o = n26269_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n26273_o = n26270_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n26275_o = write_in ? n26267_o : n26273_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n26277_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n26280_o = n26277_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n26302_o = write_in ? n26261_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n26258_o)
    if (n26258_o)
      n26303_q <= 8'b00000000;
    else
      n26303_q <= n26302_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n26258_o)
    if (n26258_o)
      n26304_q <= 8'b00000000;
    else
      n26304_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n26258_o)
    if (n26258_o)
      n26305_q <= 8'b00000000;
    else
      n26305_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n26258_o)
    if (n26258_o)
      n26307_q <= 1'b0;
    else
      n26307_q <= n26280_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n26258_o)
    if (n26258_o)
      n26308_q <= 1'b0;
    else
      n26308_q <= n26275_o;
endmodule

module ramw2_16_16_4_4_776_776
  (input  clock,
   input  clock_x2,
   input  [3:0] address_a,
   input  [775:0] data_a,
   input  wren_a,
   input  [3:0] address_b,
   output [775:0] q_b);
  wire [387:0] data;
  wire [387:0] data_r;
  wire [4:0] waddress;
  wire [3:0] waddress_r;
  wire [4:0] raddress;
  wire [3:0] raddress_r;
  wire [387:0] q;
  wire [387:0] q_latch;
  wire wren;
  wire wren_r;
  wire [387:0] n26201_o;
  wire n26202_o;
  wire [387:0] n26203_o;
  wire n26204_o;
  wire [3:0] n26205_o;
  wire n26206_o;
  wire n26207_o;
  wire [3:0] n26208_o;
  wire n26209_o;
  wire n26210_o;
  wire n26211_o;
  wire n26212_o;
  wire n26213_o;
  wire [387:0] sync_latch_i_n26214;
  wire [387:0] sync_latch_i_data_out;
  wire [387:0] n26220_o;
  wire [387:0] ram_i_n26226;
  wire [387:0] ram_i_q_b;
  reg [387:0] n26229_q;
  wire [4:0] n26230_o;
  reg [3:0] n26231_q;
  wire [4:0] n26232_o;
  reg [3:0] n26233_q;
  reg n26234_q;
  wire [775:0] n26235_o;
  assign q_b = n26235_o;
  /* ../../HW/src/util/ramw2.vhd:54:8  */
  assign data = n26203_o; // (signal)
  /* ../../HW/src/util/ramw2.vhd:55:8  */
  assign data_r = n26229_q; // (signal)
  /* ../../HW/src/util/ramw2.vhd:56:8  */
  assign waddress = n26230_o; // (signal)
  /* ../../HW/src/util/ramw2.vhd:57:8  */
  assign waddress_r = n26231_q; // (signal)
  /* ../../HW/src/util/ramw2.vhd:58:8  */
  assign raddress = n26232_o; // (signal)
  /* ../../HW/src/util/ramw2.vhd:59:8  */
  assign raddress_r = n26233_q; // (signal)
  /* ../../HW/src/util/ramw2.vhd:60:8  */
  assign q = ram_i_n26226; // (signal)
  /* ../../HW/src/util/ramw2.vhd:61:8  */
  assign q_latch = sync_latch_i_n26214; // (signal)
  /* ../../HW/src/util/ramw2.vhd:62:8  */
  assign wren = n26213_o; // (signal)
  /* ../../HW/src/util/ramw2.vhd:63:8  */
  assign wren_r = n26234_q; // (signal)
  /* ../../HW/src/util/ramw2.vhd:66:15  */
  assign n26201_o = data_a[775:388];
  /* ../../HW/src/util/ramw2.vhd:66:66  */
  assign n26202_o = ~clock;
  /* ../../HW/src/util/ramw2.vhd:66:56  */
  assign n26203_o = n26202_o ? n26201_o : data_r;
  /* ../../HW/src/util/ramw2.vhd:67:61  */
  assign n26204_o = ~clock;
  /* ../../HW/src/util/ramw2.vhd:67:51  */
  assign n26205_o = n26204_o ? address_a : waddress_r;
  /* ../../HW/src/util/ramw2.vhd:68:17  */
  assign n26206_o = ~clock;
  /* ../../HW/src/util/ramw2.vhd:69:61  */
  assign n26207_o = ~clock;
  /* ../../HW/src/util/ramw2.vhd:69:51  */
  assign n26208_o = n26207_o ? address_b : raddress_r;
  /* ../../HW/src/util/ramw2.vhd:70:17  */
  assign n26209_o = ~clock;
  /* ../../HW/src/util/ramw2.vhd:73:17  */
  assign n26210_o = wren_r & clock;
  /* ../../HW/src/util/ramw2.vhd:73:44  */
  assign n26211_o = ~clock;
  /* ../../HW/src/util/ramw2.vhd:73:39  */
  assign n26212_o = wren_a & n26211_o;
  /* ../../HW/src/util/ramw2.vhd:73:28  */
  assign n26213_o = n26210_o | n26212_o;
  /* ../../HW/src/util/ramw2.vhd:84:17  */
  assign sync_latch_i_n26214 = sync_latch_i_data_out; // (signal)
  /* ../../HW/src/util/ramw2.vhd:75:1  */
  sync_latch_388 sync_latch_i (
    .enable_in(clock),
    .data_in(q),
    .data_out(sync_latch_i_data_out));
  /* ../../HW/src/util/ramw2.vhd:90:23  */
  assign n26220_o = data_a[387:0];
  /* ../../HW/src/util/ramw2.vhd:110:14  */
  assign ram_i_n26226 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/ramw2.vhd:97:1  */
  dpram_32_32_5_5_388_388 ram_i (
    .address_a(waddress),
    .clock(clock_x2),
    .data_a(data),
    .wren_a(wren),
    .address_b(raddress),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  always @(posedge clock)
    n26229_q <= n26220_o;
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  assign n26230_o = {n26205_o, n26206_o};
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  always @(posedge clock)
    n26231_q <= address_a;
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  assign n26232_o = {n26208_o, n26209_o};
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  always @(posedge clock)
    n26233_q <= address_b;
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  always @(posedge clock)
    n26234_q <= wren_a;
  /* ../../HW/src/util/ramw2.vhd:89:4  */
  assign n26235_o = {q_latch, q};
endmodule

module dp_fifo
  (input  clock_in,
   input  reset_in,
   input  [1517:0] writedata_in,
   input  wreq_in,
   input  rdreq1_in,
   input  rdreq2_in,
   output [1517:0] readdata1_out,
   output [1517:0] readdata2_out,
   output valid1_out,
   output valid2_out,
   output full_out,
   output [7:0] fifo_avail_out);
  wire [7:0] fifo_avail_r;
  wire [7:0] wrusedw;
  wire full_r;
  wire empty;
  wire empty_normal;
  wire [1517:0] readdata;
  wire [1517:0] readdata_normal;
  wire wreq_normal;
  wire rdreq;
  wire rdreq_normal;
  wire valid1;
  wire valid2;
  wire [1517:0] readdata1;
  wire [1517:0] readdata2;
  wire valid1_r;
  wire valid2_r;
  wire [1517:0] readdata1_r;
  wire [1517:0] readdata2_r;
  wire rdreq1_r;
  wire rdreq2_r;
  wire writeready;
  wire pause;
  wire readdata1_valid_r;
  wire readdata2_valid_r;
  wire n26050_o;
  wire n26051_o;
  wire gen1_fifo_i_n26052;
  wire [1517:0] gen1_fifo_i_n26053;
  wire gen1_fifo_i_n26054;
  wire [7:0] gen1_fifo_i_n26055;
  wire gen1_fifo_i_writeready_out;
  wire [1517:0] gen1_fifo_i_q_out;
  wire gen1_fifo_i_empty_out;
  wire [7:0] gen1_fifo_i_wused_out;
  wire n26065_o;
  wire n26066_o;
  wire n26067_o;
  wire n26069_o;
  wire n26072_o;
  wire n26074_o;
  wire n26075_o;
  wire n26076_o;
  wire n26077_o;
  wire n26078_o;
  wire n26079_o;
  wire n26080_o;
  wire n26081_o;
  wire n26082_o;
  wire n26083_o;
  wire n26084_o;
  wire n26085_o;
  wire n26116_o;
  wire n26117_o;
  wire n26118_o;
  wire n26119_o;
  wire n26120_o;
  wire n26122_o;
  wire n26123_o;
  wire [1517:0] n26124_o;
  wire n26125_o;
  wire n26127_o;
  wire n26128_o;
  wire [1517:0] n26129_o;
  wire [1517:0] n26130_o;
  wire n26131_o;
  wire n26132_o;
  wire n26133_o;
  wire n26134_o;
  wire n26135_o;
  wire n26136_o;
  wire n26137_o;
  wire n26139_o;
  wire n26140_o;
  wire n26141_o;
  wire n26142_o;
  wire n26143_o;
  wire n26144_o;
  wire n26145_o;
  wire n26146_o;
  wire n26147_o;
  wire n26150_o;
  wire n26151_o;
  wire [1517:0] n26152_o;
  wire n26153_o;
  wire n26154_o;
  wire n26155_o;
  wire n26157_o;
  wire n26158_o;
  wire [1517:0] n26159_o;
  wire n26160_o;
  wire n26161_o;
  wire n26162_o;
  wire [1517:0] n26163_o;
  wire n26164_o;
  wire n26166_o;
  wire n26167_o;
  wire [1517:0] n26168_o;
  wire [1517:0] n26169_o;
  wire n26173_o;
  wire [7:0] n26175_o;
  wire [7:0] n26176_o;
  wire n26178_o;
  wire n26181_o;
  reg [7:0] n26189_q;
  reg n26190_q;
  reg n26191_q;
  reg n26192_q;
  reg [1517:0] n26193_q;
  reg [1517:0] n26194_q;
  reg n26195_q;
  reg n26196_q;
  reg n26198_q;
  reg n26199_q;
  assign readdata1_out = readdata1_r;
  assign readdata2_out = readdata2_r;
  assign valid1_out = readdata1_valid_r;
  assign valid2_out = readdata2_valid_r;
  assign full_out = n26051_o;
  assign fifo_avail_out = fifo_avail_r;
  /* ../../HW/src/dp/dp_fifo.vhd:56:8  */
  assign fifo_avail_r = n26189_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:57:8  */
  assign wrusedw = gen1_fifo_i_n26055; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:58:8  */
  assign full_r = n26190_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:59:8  */
  assign empty = empty_normal; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:60:8  */
  assign empty_normal = gen1_fifo_i_n26054; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:215:1  */
  assign readdata = readdata_normal; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:62:8  */
  assign readdata_normal = gen1_fifo_i_n26053; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:63:8  */
  assign wreq_normal = wreq_in; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:64:8  */
  assign rdreq = n26164_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:65:8  */
  assign rdreq_normal = n26067_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:66:8  */
  assign valid1 = n26166_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:67:8  */
  assign valid2 = n26167_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:68:8  */
  assign readdata1 = n26168_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:69:8  */
  assign readdata2 = n26169_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:70:8  */
  assign valid1_r = n26191_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:71:8  */
  assign valid2_r = n26192_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:72:8  */
  assign readdata1_r = n26193_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:73:8  */
  assign readdata2_r = n26194_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:74:8  */
  assign rdreq1_r = n26195_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:75:8  */
  assign rdreq2_r = n26196_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:77:8  */
  assign writeready = gen1_fifo_i_n26052; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:78:8  */
  assign pause = n26069_o; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:79:8  */
  assign readdata1_valid_r = n26198_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:80:8  */
  assign readdata2_valid_r = n26199_q; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:86:24  */
  assign n26050_o = ~writeready;
  /* ../../HW/src/dp/dp_fifo.vhd:86:20  */
  assign n26051_o = full_r | n26050_o;
  /* ../../HW/src/dp/dp_fifo.vhd:102:25  */
  assign gen1_fifo_i_n26052 = gen1_fifo_i_writeready_out; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:104:16  */
  assign gen1_fifo_i_n26053 = gen1_fifo_i_q_out; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:106:20  */
  assign gen1_fifo_i_n26054 = gen1_fifo_i_empty_out; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:105:20  */
  assign gen1_fifo_i_n26055 = gen1_fifo_i_wused_out; // (signal)
  /* ../../HW/src/dp/dp_fifo.vhd:90:1  */
  scfifow_1518_8 gen1_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(writedata_in),
    .write_in(wreq_normal),
    .read_in(rdreq_normal),
    .writeready_out(gen1_fifo_i_writeready_out),
    .q_out(gen1_fifo_i_q_out),
    .empty_out(gen1_fifo_i_empty_out),
    .wused_out(gen1_fifo_i_wused_out));
  /* ../../HW/src/dp/dp_fifo.vhd:148:52  */
  assign n26065_o = ~empty_normal;
  /* ../../HW/src/dp/dp_fifo.vhd:148:36  */
  assign n26066_o = n26065_o & rdreq;
  /* ../../HW/src/dp/dp_fifo.vhd:148:21  */
  assign n26067_o = n26066_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fifo.vhd:154:20  */
  assign n26069_o = rdreq1_in | rdreq2_in;
  /* ../../HW/src/dp/dp_fifo.vhd:158:16  */
  assign n26072_o = ~reset_in;
  /* ../../HW/src/dp/dp_fifo.vhd:177:45  */
  assign n26074_o = ~pause;
  /* ../../HW/src/dp/dp_fifo.vhd:177:40  */
  assign n26075_o = valid1 & n26074_o;
  /* ../../HW/src/dp/dp_fifo.vhd:177:66  */
  assign n26076_o = ~valid1;
  /* ../../HW/src/dp/dp_fifo.vhd:177:78  */
  assign n26077_o = n26076_o & valid2;
  /* ../../HW/src/dp/dp_fifo.vhd:177:61  */
  assign n26078_o = ~n26077_o;
  /* ../../HW/src/dp/dp_fifo.vhd:177:56  */
  assign n26079_o = n26075_o & n26078_o;
  /* ../../HW/src/dp/dp_fifo.vhd:178:45  */
  assign n26080_o = ~pause;
  /* ../../HW/src/dp/dp_fifo.vhd:178:40  */
  assign n26081_o = valid2 & n26080_o;
  /* ../../HW/src/dp/dp_fifo.vhd:178:66  */
  assign n26082_o = ~valid1;
  /* ../../HW/src/dp/dp_fifo.vhd:178:78  */
  assign n26083_o = n26082_o & valid2;
  /* ../../HW/src/dp/dp_fifo.vhd:178:61  */
  assign n26084_o = ~n26083_o;
  /* ../../HW/src/dp/dp_fifo.vhd:178:56  */
  assign n26085_o = n26081_o & n26084_o;
  /* ../../HW/src/dp/dp_fifo.vhd:198:17  */
  assign n26116_o = valid2_r & valid1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:205:17  */
  assign n26117_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:208:16  */
  assign n26118_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:211:17  */
  assign n26119_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:213:16  */
  assign n26120_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:209:4  */
  assign n26122_o = rdreq2_r ? n26120_o : 1'b0;
  /* ../../HW/src/dp/dp_fifo.vhd:209:4  */
  assign n26123_o = rdreq2_r ? n26119_o : valid2_r;
  /* ../../HW/src/dp/dp_fifo.vhd:209:4  */
  assign n26124_o = rdreq2_r ? readdata : readdata2_r;
  /* ../../HW/src/dp/dp_fifo.vhd:200:4  */
  assign n26125_o = rdreq1_r ? n26118_o : n26122_o;
  /* ../../HW/src/dp/dp_fifo.vhd:200:4  */
  assign n26127_o = rdreq1_r ? 1'b1 : valid1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:200:4  */
  assign n26128_o = rdreq1_r ? n26117_o : n26123_o;
  /* ../../HW/src/dp/dp_fifo.vhd:200:4  */
  assign n26129_o = rdreq1_r ? readdata2_r : readdata1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:200:4  */
  assign n26130_o = rdreq1_r ? readdata : n26124_o;
  /* ../../HW/src/dp/dp_fifo.vhd:215:32  */
  assign n26131_o = ~valid2_r;
  /* ../../HW/src/dp/dp_fifo.vhd:215:20  */
  assign n26132_o = n26131_o & valid1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:219:17  */
  assign n26133_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:221:16  */
  assign n26134_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:223:17  */
  assign n26135_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:225:16  */
  assign n26136_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:217:4  */
  assign n26137_o = rdreq1_r ? n26134_o : n26136_o;
  /* ../../HW/src/dp/dp_fifo.vhd:217:4  */
  assign n26139_o = rdreq1_r ? 1'b0 : valid1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:217:4  */
  assign n26140_o = rdreq1_r ? n26133_o : n26135_o;
  /* ../../HW/src/dp/dp_fifo.vhd:227:15  */
  assign n26141_o = ~valid1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:227:20  */
  assign n26142_o = valid2_r & n26141_o;
  /* ../../HW/src/dp/dp_fifo.vhd:230:17  */
  assign n26143_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:232:16  */
  assign n26144_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:237:17  */
  assign n26145_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:239:16  */
  assign n26146_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:229:4  */
  assign n26147_o = rdreq2_r ? n26144_o : n26146_o;
  /* ../../HW/src/dp/dp_fifo.vhd:229:4  */
  assign n26150_o = rdreq2_r ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fifo.vhd:229:4  */
  assign n26151_o = rdreq2_r ? n26143_o : n26145_o;
  /* ../../HW/src/dp/dp_fifo.vhd:229:4  */
  assign n26152_o = rdreq2_r ? readdata1_r : readdata2_r;
  /* ../../HW/src/dp/dp_fifo.vhd:243:14  */
  assign n26153_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:245:13  */
  assign n26154_o = ~empty;
  /* ../../HW/src/dp/dp_fifo.vhd:227:1  */
  assign n26155_o = n26142_o ? n26147_o : n26154_o;
  /* ../../HW/src/dp/dp_fifo.vhd:227:1  */
  assign n26157_o = n26142_o ? n26150_o : 1'b0;
  /* ../../HW/src/dp/dp_fifo.vhd:227:1  */
  assign n26158_o = n26142_o ? n26151_o : n26153_o;
  /* ../../HW/src/dp/dp_fifo.vhd:227:1  */
  assign n26159_o = n26142_o ? n26152_o : readdata1_r;
  /* ../../HW/src/dp/dp_fifo.vhd:215:1  */
  assign n26160_o = n26132_o ? n26137_o : n26155_o;
  /* ../../HW/src/dp/dp_fifo.vhd:215:1  */
  assign n26161_o = n26132_o ? n26139_o : n26157_o;
  /* ../../HW/src/dp/dp_fifo.vhd:215:1  */
  assign n26162_o = n26132_o ? n26140_o : n26158_o;
  /* ../../HW/src/dp/dp_fifo.vhd:215:1  */
  assign n26163_o = n26132_o ? readdata1_r : n26159_o;
  /* ../../HW/src/dp/dp_fifo.vhd:198:1  */
  assign n26164_o = n26116_o ? n26125_o : n26160_o;
  /* ../../HW/src/dp/dp_fifo.vhd:198:1  */
  assign n26166_o = n26116_o ? n26127_o : n26161_o;
  /* ../../HW/src/dp/dp_fifo.vhd:198:1  */
  assign n26167_o = n26116_o ? n26128_o : n26162_o;
  /* ../../HW/src/dp/dp_fifo.vhd:198:1  */
  assign n26168_o = n26116_o ? n26129_o : n26163_o;
  /* ../../HW/src/dp/dp_fifo.vhd:198:1  */
  assign n26169_o = n26116_o ? n26130_o : readdata;
  /* ../../HW/src/dp/dp_fifo.vhd:253:16  */
  assign n26173_o = ~reset_in;
  /* ../../HW/src/dp/dp_fifo.vhd:258:30  */
  assign n26175_o = ~wrusedw;
  /* ../../HW/src/dp/dp_fifo.vhd:259:25  */
  assign n26176_o = ~wrusedw;
  /* ../../HW/src/dp/dp_fifo.vhd:259:38  */
  assign n26178_o = $unsigned(n26176_o) < $unsigned(8'b00000100);
  /* ../../HW/src/dp/dp_fifo.vhd:259:13  */
  assign n26181_o = n26178_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fifo.vhd:257:9  */
  always @(posedge clock_in or posedge n26173_o)
    if (n26173_o)
      n26189_q <= 8'b00000000;
    else
      n26189_q <= n26175_o;
  /* ../../HW/src/dp/dp_fifo.vhd:257:9  */
  always @(posedge clock_in or posedge n26173_o)
    if (n26173_o)
      n26190_q <= 1'b0;
    else
      n26190_q <= n26181_o;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26191_q <= 1'b0;
    else
      n26191_q <= valid1;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26192_q <= 1'b0;
    else
      n26192_q <= valid2;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26193_q <= 1518'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n26193_q <= readdata1;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26194_q <= 1518'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n26194_q <= readdata2;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26195_q <= 1'b0;
    else
      n26195_q <= rdreq1_in;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26196_q <= 1'b0;
    else
      n26196_q <= rdreq2_in;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26198_q <= 1'b0;
    else
      n26198_q <= n26079_o;
  /* ../../HW/src/dp/dp_fifo.vhd:169:9  */
  always @(posedge clock_in or posedge n26072_o)
    if (n26072_o)
      n26199_q <= 1'b0;
    else
      n26199_q <= n26085_o;
endmodule

module scfifo_64_8_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [63:0] data_in,
   input  write_in,
   input  read_in,
   output [63:0] q_out,
   output [7:0] ravail_out,
   output [7:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [63:0] q;
  wire [7:0] address_a;
  wire [7:0] address_b;
  wire [7:0] waddr_r;
  wire [7:0] waddr_rr;
  wire [7:0] raddr_r;
  wire [7:0] raddr;
  wire [7:0] ravail;
  wire [7:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [63:0] ram_i_n25977;
  wire [63:0] ram_i_q_b;
  wire [7:0] n25980_o;
  wire [7:0] n25981_o;
  wire n25982_o;
  wire n25985_o;
  wire n25986_o;
  wire [7:0] n25989_o;
  wire [7:0] n25990_o;
  wire n25993_o;
  wire [7:0] n25996_o;
  wire [7:0] n25998_o;
  wire n25999_o;
  wire n26002_o;
  wire [7:0] n26004_o;
  wire n26005_o;
  wire n26008_o;
  wire n26010_o;
  wire n26012_o;
  wire n26015_o;
  wire [7:0] n26037_o;
  reg [7:0] n26038_q;
  reg [7:0] n26039_q;
  reg [7:0] n26040_q;
  reg n26042_q;
  reg n26043_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n25982_o;
  assign full_out = full_r;
  assign almost_full_out = n25986_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n25977; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n26038_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n26039_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n26040_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n25990_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n25980_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n25981_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n26042_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n26043_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n25977 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_256_256_8_8_64_64 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n25980_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n25981_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n25982_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n25985_o = $unsigned(wused) >= $unsigned(8'b00000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n25986_o = n25985_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n25989_o = raddr_r + 8'b00000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n25990_o = read_in ? n25989_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n25993_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n25996_o = waddr_r + 8'b00000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n25998_o = waddr_r + 8'b00000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n25999_o = n25998_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n26002_o = n25999_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n26004_o = waddr_r + 8'b00000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n26005_o = n26004_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n26008_o = n26005_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n26010_o = write_in ? n26002_o : n26008_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n26012_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n26015_o = n26012_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n26037_o = write_in ? n25996_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n25993_o)
    if (n25993_o)
      n26038_q <= 8'b00000000;
    else
      n26038_q <= n26037_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n25993_o)
    if (n25993_o)
      n26039_q <= 8'b00000000;
    else
      n26039_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n25993_o)
    if (n25993_o)
      n26040_q <= 8'b00000000;
    else
      n26040_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n25993_o)
    if (n25993_o)
      n26042_q <= 1'b0;
    else
      n26042_q <= n26015_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n25993_o)
    if (n25993_o)
      n26043_q <= 1'b0;
    else
      n26043_q <= n26010_o;
endmodule

module pcore_1_3
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire dp_wr_fork;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire dp_wr_fork_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n24802_o;
  wire n24803_o;
  wire n24804_o;
  wire n24807_o;
  wire [4:0] n24895_o;
  wire n24896_o;
  wire [4:0] n24897_o;
  wire n24898_o;
  wire [2:0] n24901_o;
  wire [4:0] n24903_o;
  wire n24904_o;
  wire n24905_o;
  wire n24906_o;
  wire n24907_o;
  wire [4:0] n24908_o;
  wire [4:0] n24909_o;
  wire [4:0] n24910_o;
  wire n24911_o;
  wire n24912_o;
  wire n24913_o;
  wire [4:0] n24914_o;
  wire n24915_o;
  wire n24916_o;
  wire [4:0] n24917_o;
  wire n24918_o;
  wire n24919_o;
  wire n24920_o;
  wire n24921_o;
  wire n24924_o;
  wire n24930_o;
  wire n24932_o;
  wire [2:0] n24934_o;
  wire n24936_o;
  wire n24937_o;
  wire n24938_o;
  wire [2:0] n24940_o;
  wire [2:0] n24942_o;
  wire [2:0] n24944_o;
  wire n24945_o;
  wire n24946_o;
  wire [21:0] n24947_o;
  wire n24948_o;
  wire [2:0] n24949_o;
  wire [1:0] n24950_o;
  wire n24951_o;
  wire [21:0] n24952_o;
  wire n24953_o;
  wire [1:0] n24954_o;
  wire [1:0] n24955_o;
  wire n24956_o;
  wire [1:0] n24957_o;
  wire [2:0] n24958_o;
  wire [2:0] n24959_o;
  wire n24964_o;
  wire n24965_o;
  wire n24966_o;
  wire n24967_o;
  wire n24968_o;
  wire n24970_o;
  wire [2:0] n24972_o;
  wire n24974_o;
  wire n24975_o;
  wire n24976_o;
  wire [2:0] n24978_o;
  wire [2:0] n24982_o;
  wire [2:0] n24984_o;
  wire n24985_o;
  wire n24986_o;
  wire [21:0] n24987_o;
  wire [5:0] n24988_o;
  wire n24989_o;
  wire [2:0] n24990_o;
  wire [1:0] n24991_o;
  wire n24992_o;
  wire [21:0] n24993_o;
  wire [2:0] n24995_o;
  wire [2:0] n24998_o;
  wire n25003_o;
  wire n25006_o;
  wire n25007_o;
  wire [21:0] n25008_o;
  wire [21:0] n25010_o;
  wire [21:0] n25011_o;
  wire [21:0] n25013_o;
  wire [21:0] n25014_o;
  wire n25016_o;
  wire n25080_o;
  wire n25149_o;
  wire n25152_o;
  wire n25153_o;
  wire [21:0] n25154_o;
  wire [21:0] n25156_o;
  wire [21:0] n25157_o;
  wire [21:0] n25159_o;
  wire [21:0] n25160_o;
  wire n25162_o;
  wire [83:0] n25163_o;
  wire [83:0] n25164_o;
  wire [83:0] n25174_o;
  wire [11:0] n25216_o;
  wire [11:0] n25217_o;
  wire n25231_o;
  wire n25233_o;
  wire [11:0] n25234_o;
  wire [11:0] n25235_o;
  wire [11:0] n25236_o;
  wire [95:0] n25238_o;
  wire [95:0] n25239_o;
  wire [1:0] n25245_o;
  wire [2:0] n25246_o;
  wire n25247_o;
  wire n25249_o;
  wire n25250_o;
  wire n25252_o;
  wire n25253_o;
  wire n25256_o;
  wire n25258_o;
  wire n25259_o;
  wire n25262_o;
  wire n25263_o;
  wire [1:0] n25265_o;
  wire [1:0] n25267_o;
  wire n25269_o;
  wire [1:0] n25271_o;
  wire [1:0] n25277_o;
  wire [2:0] n25278_o;
  wire [4:0] n25279_o;
  wire n25282_o;
  wire [95:0] n25283_o;
  wire [95:0] n25285_o;
  wire n25287_o;
  wire n25292_o;
  wire n25343_o;
  wire n25346_o;
  wire [2:0] n25347_o;
  wire [11:0] n25348_o;
  wire n25350_o;
  wire [11:0] n25351_o;
  wire n25353_o;
  wire [11:0] n25354_o;
  wire n25356_o;
  wire [11:0] n25357_o;
  wire n25359_o;
  wire [11:0] n25360_o;
  wire n25362_o;
  wire [11:0] n25363_o;
  wire n25365_o;
  wire [11:0] n25366_o;
  wire n25368_o;
  wire [11:0] n25369_o;
  wire [6:0] n25370_o;
  wire [11:0] n25371_o;
  reg [11:0] n25372_o;
  wire [11:0] n25373_o;
  reg [11:0] n25374_o;
  wire [11:0] n25375_o;
  reg [11:0] n25376_o;
  wire [11:0] n25377_o;
  reg [11:0] n25378_o;
  wire [11:0] n25379_o;
  reg [11:0] n25380_o;
  wire [11:0] n25381_o;
  reg [11:0] n25382_o;
  wire [11:0] n25383_o;
  reg [11:0] n25384_o;
  wire [11:0] n25385_o;
  reg [11:0] n25386_o;
  wire n25388_o;
  wire n25391_o;
  wire [95:0] n25392_o;
  wire [95:0] n25393_o;
  wire [95:0] n25394_o;
  wire [95:0] n25395_o;
  wire [95:0] n25396_o;
  wire n25398_o;
  wire [2:0] n25400_o;
  wire [2:0] n25402_o;
  wire n25407_o;
  wire [12:0] xregister_file_i_n25456;
  wire [255:0] xregister_file_i_n25457;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n25462;
  wire [12:0] iregister_i_n25463;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n25470_o;
  wire n25472_o;
  wire n25473_o;
  wire n25475_o;
  wire n25476_o;
  wire n25479_o;
  wire n25481_o;
  wire n25482_o;
  wire n25485_o;
  wire n25486_o;
  wire [4:0] n25494_o;
  wire n25495_o;
  wire [4:0] n25496_o;
  wire [4:0] n25499_o;
  wire [4:0] n25500_o;
  wire [4:0] n25501_o;
  wire n25502_o;
  wire n25503_o;
  wire n25504_o;
  wire n25505_o;
  wire n25506_o;
  wire n25507_o;
  wire n25508_o;
  wire n25509_o;
  wire n25510_o;
  wire n25513_o;
  wire [31:0] n25515_o;
  wire [11:0] n25516_o;
  wire [11:0] n25517_o;
  wire [31:0] alu_0_i_n25518;
  wire alu_0_i_n25519;
  wire [11:0] alu_0_i_n25520;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n25527_o;
  wire [11:0] n25528_o;
  wire [11:0] n25529_o;
  wire [31:0] alu_1_i_n25530;
  wire alu_1_i_n25531;
  wire [11:0] alu_1_i_n25532;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n25539_o;
  wire [11:0] n25540_o;
  wire [11:0] n25541_o;
  wire [31:0] alu_2_i_n25542;
  wire alu_2_i_n25543;
  wire [11:0] alu_2_i_n25544;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n25551_o;
  wire [11:0] n25552_o;
  wire [11:0] n25553_o;
  wire [31:0] alu_3_i_n25554;
  wire alu_3_i_n25555;
  wire [11:0] alu_3_i_n25556;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n25563_o;
  wire [11:0] n25564_o;
  wire [11:0] n25565_o;
  wire [31:0] alu_4_i_n25566;
  wire alu_4_i_n25567;
  wire [11:0] alu_4_i_n25568;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n25575_o;
  wire [11:0] n25576_o;
  wire [11:0] n25577_o;
  wire [31:0] alu_5_i_n25578;
  wire alu_5_i_n25579;
  wire [11:0] alu_5_i_n25580;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n25587_o;
  wire [11:0] n25588_o;
  wire [11:0] n25589_o;
  wire [31:0] alu_6_i_n25590;
  wire alu_6_i_n25591;
  wire [11:0] alu_6_i_n25592;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n25599_o;
  wire [11:0] n25600_o;
  wire [11:0] n25601_o;
  wire [31:0] alu_7_i_n25602;
  wire alu_7_i_n25603;
  wire [11:0] alu_7_i_n25604;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n25611_o;
  wire n25612_o;
  wire [12:0] ialu_i_n25613;
  wire ialu_i_n25614;
  wire ialu_i_n25615;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n25624;
  wire [95:0] register_bank_i_n25625;
  wire [16:0] n25626_o;
  wire [16:0] n25627_o;
  wire [95:0] register_bank_i_n25628;
  wire register_bank_i_n25629;
  wire register_bank_i_n25630;
  wire [2:0] register_bank_i_n25631;
  wire [2:0] register_bank_i_n25632;
  wire [1:0] register_bank_i_n25633;
  wire [2:0] register_bank_i_n25634;
  wire [2:0] register_bank_i_n25635;
  wire register_bank_i_n25636;
  wire [1:0] register_bank_i_n25637;
  wire [1:0] register_bank_i_n25638;
  wire register_bank_i_n25639;
  wire [1:0] register_bank_i_n25640;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n25673;
  wire instr_decoder2_i_n25674;
  wire [3:0] instr_decoder2_i_n25675;
  wire instr_decoder2_i_n25676;
  wire instr_decoder2_i_n25677;
  wire instr_decoder2_i_n25678;
  wire instr_decoder2_i_n25679;
  wire [11:0] instr_decoder2_i_n25680;
  wire [11:0] instr_decoder2_i_n25681;
  wire [11:0] instr_decoder2_i_n25682;
  wire instr_decoder2_i_n25683;
  wire instr_decoder2_i_n25684;
  wire instr_decoder2_i_n25685;
  wire [7:0] instr_decoder2_i_n25686;
  wire instr_decoder2_i_n25687;
  wire [11:0] instr_decoder2_i_n25688;
  wire instr_decoder2_i_n25689;
  wire instr_decoder2_i_n25690;
  wire [3:0] instr_decoder2_i_n25691;
  wire [3:0] instr_decoder2_i_n25692;
  wire instr_decoder2_i_n25693;
  wire instr_decoder2_i_n25694;
  wire [2:0] instr_decoder2_i_n25695;
  wire [12:0] instr_decoder2_i_n25696;
  wire instr_decoder2_i_n25697;
  wire [4:0] instr_decoder2_i_n25698;
  wire [12:0] instr_decoder2_i_n25699;
  wire [12:0] instr_decoder2_i_n25700;
  wire [7:0] instr_decoder2_i_n25701;
  wire [7:0] instr_decoder2_i_n25702;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n25763;
  wire instr_dispatch2_i1_n25764;
  wire [11:0] instr_dispatch2_i1_n25765;
  wire [11:0] instr_dispatch2_i1_n25766;
  wire instr_dispatch2_i1_n25767;
  wire instr_dispatch2_i1_n25768;
  wire instr_dispatch2_i1_n25769;
  wire instr_dispatch2_i1_n25770;
  wire instr_dispatch2_i1_n25771;
  wire instr_dispatch2_i1_n25772;
  wire instr_dispatch2_i1_n25773;
  wire instr_dispatch2_i1_n25774;
  wire [11:0] instr_dispatch2_i1_n25775;
  wire [7:0] instr_dispatch2_i1_n25776;
  wire [95:0] instr_dispatch2_i1_n25777;
  wire [7:0] instr_dispatch2_i1_n25778;
  wire [95:0] instr_dispatch2_i1_n25779;
  wire [95:0] instr_dispatch2_i1_n25780;
  wire [11:0] instr_dispatch2_i1_n25781;
  wire [4:0] instr_dispatch2_i1_n25782;
  wire [3:0] instr_dispatch2_i1_n25783;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n25829_o;
  wire [95:0] n25830_o;
  wire [7:0] n25831_o;
  wire [95:0] n25832_o;
  reg [95:0] n25833_q;
  wire [95:0] n25834_o;
  reg [95:0] n25835_q;
  reg n25836_q;
  reg n25837_q;
  wire n25838_o;
  reg n25839_q;
  wire [1:0] n25840_o;
  reg [1:0] n25841_q;
  wire [1:0] n25842_o;
  reg [1:0] n25843_q;
  wire [2:0] n25844_o;
  reg [2:0] n25845_q;
  wire [2:0] n25846_o;
  reg [2:0] n25847_q;
  wire n25848_o;
  reg n25849_q;
  wire [1:0] n25850_o;
  reg [1:0] n25851_q;
  reg [2:0] n25852_q;
  reg [2:0] n25853_q;
  reg [1:0] n25854_q;
  reg [2:0] n25857_q;
  reg [2:0] n25858_q;
  reg n25859_q;
  reg [1:0] n25860_q;
  reg [1:0] n25861_q;
  reg n25862_q;
  reg [1:0] n25863_q;
  reg [21:0] n25864_q;
  reg [2:0] n25865_q;
  reg [21:0] n25866_q;
  reg [95:0] n25867_q;
  wire n25868_o;
  reg n25869_q;
  wire n25870_o;
  reg n25871_q;
  wire n25872_o;
  reg n25873_q;
  wire n25874_o;
  reg n25875_q;
  reg [21:0] n25876_q;
  reg [21:0] n25877_q;
  wire [5:0] n25878_o;
  reg [5:0] n25879_q;
  wire n25880_o;
  reg n25881_q;
  wire [2:0] n25884_o;
  reg [2:0] n25885_q;
  wire [1:0] n25886_o;
  reg [1:0] n25887_q;
  wire n25888_o;
  reg n25889_q;
  wire [21:0] n25890_o;
  reg [21:0] n25891_q;
  wire n25892_o;
  reg n25893_q;
  wire [2:0] n25894_o;
  reg [2:0] n25895_q;
  wire [1:0] n25896_o;
  reg [1:0] n25897_q;
  wire n25898_o;
  wire n25899_o;
  wire n25900_o;
  reg n25901_q;
  wire n25902_o;
  wire n25903_o;
  wire [21:0] n25904_o;
  reg [21:0] n25905_q;
  wire n25906_o;
  reg n25907_q;
  wire [1:0] n25908_o;
  reg [1:0] n25909_q;
  wire [1:0] n25910_o;
  reg [1:0] n25911_q;
  wire n25912_o;
  reg n25913_q;
  wire [1:0] n25914_o;
  reg [1:0] n25915_q;
  reg [83:0] n25916_q;
  wire [95:0] n25917_o;
  reg [2:0] n25918_q;
  reg [2:0] n25919_q;
  reg [2:0] n25920_q;
  reg [79:0] n25922_q;
  reg [31:0] n25923_q;
  reg n25924_q;
  reg n25925_q;
  reg n25926_q;
  reg [1:0] n25927_q;
  reg [3:0] n25928_q;
  reg n25929_q;
  reg [3:0] n25930_q;
  reg n25931_q;
  reg [3:0] n25932_q;
  reg n25933_q;
  reg n25934_q;
  reg [1:0] n25935_q;
  reg [27:0] n25936_q;
  reg n25937_q;
  reg n25938_q;
  reg n25940_q;
  reg n25941_q;
  reg n25943_q;
  reg n25944_q;
  reg n25945_q;
  reg [21:0] n25946_q;
  reg n25947_q;
  reg [21:0] n25948_q;
  reg [21:0] n25949_q;
  reg n25950_q;
  reg [21:0] n25951_q;
  reg [5:0] n25952_q;
  reg n25953_q;
  reg n25954_q;
  reg n25955_q;
  reg [2:0] n25956_q;
  reg [1:0] n25957_q;
  reg n25958_q;
  reg n25959_q;
  reg [2:0] n25960_q;
  reg [1:0] n25961_q;
  reg n25962_q;
  reg [1:0] n25963_q;
  reg [1:0] n25964_q;
  reg n25965_q;
  reg [1:0] n25966_q;
  reg [95:0] n25967_q;
  reg n25968_q;
  wire [2:0] n25969_o;
  wire [2:0] n25970_o;
  assign i_y_neg_out = n25611_o;
  assign i_y_zero_out = n25612_o;
  assign dp_readdata_out = n25285_o;
  assign dp_readdata_vm_out = n25287_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n25969_o;
  assign dp_read_vaddr_out = n25970_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n25265_o;
  assign dp_read_data_type_out = n25267_o;
  assign dp_read_stream_out = n25269_o;
  assign dp_read_stream_id_out = n25271_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n25624; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n25625; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n25763; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n25764; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n25772; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n25769; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n25770; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n25771; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n25777; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n25778; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n25680; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n25681; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n25682; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n25463; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n25697; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n25673; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n25779; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n25780; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n25781; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n25829_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n25830_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n25831_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n25782; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n25783; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n25675; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n25513_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n25486_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n25279_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n25765; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n25766; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n25775; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n25776; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n25277_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n25278_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n25674; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n25679; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n25676; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n25677; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n25678; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n25687; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n25688; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n25683; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n25684; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n25685; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n25686; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n25767; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n25768; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n25774; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n25689; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n25690; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n25691; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n25462; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n25692; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n25693; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n25694; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n25695; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n25696; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n25833_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n25835_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n25836_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n25837_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n25839_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n25841_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n25843_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n25845_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n25847_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n25849_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n25851_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n25698; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n25699; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n25700; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n25613; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n25614; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n25615; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n25773; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n25701; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n25702; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n25456; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n25457; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n24945_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n24946_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n24985_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:191:8  */
  assign dp_wr_fork = n24986_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n24947_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n24987_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n24988_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n24989_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n24990_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n24991_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n24992_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n24993_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n24948_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n24949_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n24950_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n24951_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n24952_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n24953_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n24954_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n24955_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n24956_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n24957_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n25239_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n24958_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n24959_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n24995_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n24998_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n25852_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n25853_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n25854_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n25857_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n25858_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n25859_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n25860_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n25861_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n25862_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n25863_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n25864_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n25865_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n25866_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n25867_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n25869_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n25871_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n25873_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:238:8  */
  assign dp_wr_fork_r = n25875_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n25876_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n25877_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n25879_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n25881_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n25885_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n25887_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n25889_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n25891_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n25893_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n25895_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n25897_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n25901_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n25905_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n25907_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n25909_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n25911_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n25913_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n25915_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n25917_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n25918_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n25919_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n25920_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n25263_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n24924_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n25630; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n25631; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n25632; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n25633; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n25634; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n25635; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n25628; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n25629; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n25636; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n25637; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n25638; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n25639; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n25640; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n24802_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n24803_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n24804_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n25922_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n25923_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n25924_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n25925_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n25926_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n25927_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n25928_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n25929_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n25930_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n25931_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n25932_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n25933_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n25934_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n25935_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n25936_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n25937_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n25938_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n25940_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n25941_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n25943_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n25944_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n25945_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n25946_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n25947_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n25948_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n25949_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n25950_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n25951_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n25952_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n25953_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n25954_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n25955_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n25956_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n25957_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n25958_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n25959_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n25960_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n25961_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n25962_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n25963_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n25964_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n25965_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n25966_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n25967_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n25968_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n24802_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n24803_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n24804_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n24807_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n24895_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n24896_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n24897_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n24898_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n24901_o = n24898_o ? 3'b001 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n24903_o = n24897_o + n24895_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n24904_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n24905_o = n24904_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n24906_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n24907_o = n24906_o & n24905_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n24908_o = n24895_o & n24897_o;
  /* ../../HW/src/pcore/pcore.vhd:104:8  */
  assign n24909_o = {n24901_o, 2'b11};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n24910_o = n24895_o & n24909_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n24911_o = n24908_o == n24910_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n24912_o = n24911_o & n24896_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n24913_o = ~n24896_o;
  /* ../../HW/src/pcore/pcore.vhd:349:1  */
  assign n24914_o = {n24901_o, 2'b11};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n24915_o = $unsigned(n24914_o) >= $unsigned(n24897_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n24916_o = n24915_o & n24913_o;
  /* ../../HW/src/pcore/pcore.vhd:349:1  */
  assign n24917_o = {n24901_o, 2'b11};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n24918_o = $unsigned(n24917_o) <= $unsigned(n24903_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n24919_o = n24918_o & n24916_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n24920_o = n24912_o | n24919_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n24921_o = n24920_o & n24907_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n24924_o = n24921_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n24930_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n24932_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n24934_o = n24932_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n24936_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n24937_o = n24936_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n24938_o = dp_read_gen_valid_in_r & n24937_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n24940_o = n24938_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n24942_o = n24938_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n24944_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24945_o = n24930_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24946_o = n24930_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24947_o = n24930_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24948_o = n24930_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24949_o = n24930_o ? n24934_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24950_o = n24930_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24951_o = n24930_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24952_o = n24930_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24953_o = n24930_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24954_o = n24930_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24955_o = n24930_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24956_o = n24930_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24957_o = n24930_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24958_o = n24930_o ? n24940_o : n24944_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n24959_o = n24930_o ? n24942_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n24964_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n24965_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n24966_o = dp_write_in_r & n24965_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n24967_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n24968_o = n24966_o & n24967_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n24970_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n24972_o = n24970_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n24974_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n24975_o = n24974_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n24976_o = dp_write_gen_valid_in_r & n24975_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n24978_o = n24976_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n24982_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n24984_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24985_o = n24964_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24986_o = n24964_o ? dp_wr_fork_in_r : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24987_o = n24964_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24988_o = n24964_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24989_o = n24964_o ? n24968_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24990_o = n24964_o ? n24972_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24991_o = n24964_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24992_o = n24964_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24993_o = n24964_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24995_o = n24964_o ? n24978_o : n24982_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n24998_o = n24964_o ? 3'b000 : n24984_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n25003_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n25006_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n25007_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n25008_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n25010_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n25011_o = n25007_o ? n25008_o : n25010_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n25013_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n25014_o = n25006_o ? n25011_o : n25013_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n25016_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n25080_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n25149_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n25152_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n25153_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n25154_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n25156_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n25157_o = n25153_o ? n25154_o : n25156_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n25159_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n25160_o = n25152_o ? n25157_o : n25159_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n25162_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n25163_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n25164_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n25174_o = n25162_o ? n25163_o : n25164_o;
  assign n25216_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n25217_o = n25149_o ? 12'b000000000000 : n25216_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n25231_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n25233_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n25234_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n25235_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n25236_o = n25233_o ? n25234_o : n25235_o;
  assign n25238_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n25236_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n25239_o = n25231_o ? n25238_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n25245_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n25246_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n25247_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n25249_o = n25245_o == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n25250_o = n25249_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n25252_o = n25246_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n25253_o = n25252_o & n25250_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n25256_o = n25253_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n25258_o = n25245_o == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n25259_o = n25258_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n25262_o = n25259_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n25263_o = n25247_o ? n25256_o : n25262_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n25265_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n25267_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n25269_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n25271_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n25277_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n25278_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n25279_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n25282_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n25283_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n25285_o = n25282_o ? 96'bZ : n25283_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n25287_o = n25282_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n25292_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n25343_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n25346_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n25347_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n25348_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n25350_o = n25347_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n25351_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n25353_o = n25347_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n25354_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n25356_o = n25347_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n25357_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n25359_o = n25347_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n25360_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n25362_o = n25347_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n25363_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n25365_o = n25347_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n25366_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n25368_o = n25347_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n25369_o = dp_readdata_vm[11:0];
  assign n25370_o = {n25368_o, n25365_o, n25362_o, n25359_o, n25356_o, n25353_o, n25350_o};
  assign n25371_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25372_o = n25371_o;
      7'b0100000: n25372_o = n25371_o;
      7'b0010000: n25372_o = n25371_o;
      7'b0001000: n25372_o = n25371_o;
      7'b0000100: n25372_o = n25371_o;
      7'b0000010: n25372_o = n25371_o;
      7'b0000001: n25372_o = n25371_o;
      default: n25372_o = n25369_o;
    endcase
  assign n25373_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25374_o = n25366_o;
      7'b0100000: n25374_o = n25373_o;
      7'b0010000: n25374_o = n25373_o;
      7'b0001000: n25374_o = n25373_o;
      7'b0000100: n25374_o = n25373_o;
      7'b0000010: n25374_o = n25373_o;
      7'b0000001: n25374_o = n25373_o;
      default: n25374_o = n25373_o;
    endcase
  assign n25375_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25376_o = n25375_o;
      7'b0100000: n25376_o = n25363_o;
      7'b0010000: n25376_o = n25375_o;
      7'b0001000: n25376_o = n25375_o;
      7'b0000100: n25376_o = n25375_o;
      7'b0000010: n25376_o = n25375_o;
      7'b0000001: n25376_o = n25375_o;
      default: n25376_o = n25375_o;
    endcase
  assign n25377_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25378_o = n25377_o;
      7'b0100000: n25378_o = n25377_o;
      7'b0010000: n25378_o = n25360_o;
      7'b0001000: n25378_o = n25377_o;
      7'b0000100: n25378_o = n25377_o;
      7'b0000010: n25378_o = n25377_o;
      7'b0000001: n25378_o = n25377_o;
      default: n25378_o = n25377_o;
    endcase
  assign n25379_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25380_o = n25379_o;
      7'b0100000: n25380_o = n25379_o;
      7'b0010000: n25380_o = n25379_o;
      7'b0001000: n25380_o = n25357_o;
      7'b0000100: n25380_o = n25379_o;
      7'b0000010: n25380_o = n25379_o;
      7'b0000001: n25380_o = n25379_o;
      default: n25380_o = n25379_o;
    endcase
  assign n25381_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25382_o = n25381_o;
      7'b0100000: n25382_o = n25381_o;
      7'b0010000: n25382_o = n25381_o;
      7'b0001000: n25382_o = n25381_o;
      7'b0000100: n25382_o = n25354_o;
      7'b0000010: n25382_o = n25381_o;
      7'b0000001: n25382_o = n25381_o;
      default: n25382_o = n25381_o;
    endcase
  assign n25383_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25384_o = n25383_o;
      7'b0100000: n25384_o = n25383_o;
      7'b0010000: n25384_o = n25383_o;
      7'b0001000: n25384_o = n25383_o;
      7'b0000100: n25384_o = n25383_o;
      7'b0000010: n25384_o = n25351_o;
      7'b0000001: n25384_o = n25383_o;
      default: n25384_o = n25383_o;
    endcase
  assign n25385_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n25370_o)
      7'b1000000: n25386_o = n25385_o;
      7'b0100000: n25386_o = n25385_o;
      7'b0010000: n25386_o = n25385_o;
      7'b0001000: n25386_o = n25385_o;
      7'b0000100: n25386_o = n25385_o;
      7'b0000010: n25386_o = n25385_o;
      7'b0000001: n25386_o = n25348_o;
      default: n25386_o = n25385_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n25388_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n25391_o = n25388_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n25392_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n25393_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n25394_o = {n25386_o, n25384_o, n25382_o, n25380_o, n25378_o, n25376_o, n25374_o, n25372_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n25395_o = n25346_o ? n25394_o : n25392_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n25396_o = n25346_o ? dp_readdata2_r : n25393_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n25398_o = n25346_o ? n25391_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n25400_o = n25346_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n25402_o = n25346_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n25407_o = dp_readena_vm ? n25398_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n25456 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n25457 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n25462 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n25463 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n25470_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n25472_o = dp_rd_pid == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n25473_o = n25472_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n25475_o = dp_rd_cid == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n25476_o = n25475_o & n25473_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n25479_o = n25476_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n25481_o = dp_rd_pid == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n25482_o = n25481_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n25485_o = n25482_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n25486_o = n25470_o ? n25479_o : n25485_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n25494_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n25495_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n25496_o = dp_mcast_addr + n25494_o;
  /* ../../HW/src/pcore/pcore.vhd:1022:1  */
  assign n25499_o = dp_wr_fork ? 5'b00011 : 5'b00111;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n25500_o = n25494_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n25501_o = n25494_o & n25499_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n25502_o = n25500_o == n25501_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n25503_o = n25502_o & n25495_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n25504_o = ~n25495_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n25505_o = $unsigned(n25499_o) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n25506_o = n25505_o & n25504_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n25507_o = $unsigned(n25499_o) <= $unsigned(n25496_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n25508_o = n25507_o & n25506_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n25509_o = n25503_o | n25508_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n25510_o = n25509_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n25513_o = n25510_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n25515_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n25516_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n25517_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n25518 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n25519 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n25520 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25515_o),
    .x1_in(n25516_o),
    .x2_in(n25517_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n25527_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n25528_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n25529_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n25530 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n25531 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n25532 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25527_o),
    .x1_in(n25528_o),
    .x2_in(n25529_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n25539_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n25540_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n25541_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n25542 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n25543 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n25544 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25539_o),
    .x1_in(n25540_o),
    .x2_in(n25541_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n25551_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n25552_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n25553_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n25554 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n25555 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n25556 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25551_o),
    .x1_in(n25552_o),
    .x2_in(n25553_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n25563_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n25564_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n25565_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n25566 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n25567 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n25568 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25563_o),
    .x1_in(n25564_o),
    .x2_in(n25565_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n25575_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n25576_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n25577_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n25578 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n25579 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n25580 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25575_o),
    .x1_in(n25576_o),
    .x2_in(n25577_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n25587_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n25588_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n25589_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n25590 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n25591 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n25592 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25587_o),
    .x1_in(n25588_o),
    .x2_in(n25589_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n25599_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n25600_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n25601_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n25602 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n25603 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n25604 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n25599_o),
    .x1_in(n25600_o),
    .x2_in(n25601_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n25611_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n25612_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n25613 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n25614 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n25615 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n25624 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n25625 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n25626_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n25627_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n25628 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n25629 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n25630 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n25631 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n25632 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n25633 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n25634 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n25635 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n25636 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n25637 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n25638 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n25639 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n25640 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n25626_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n25627_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n25673 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n25674 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n25675 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n25676 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n25677 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n25678 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n25679 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n25680 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n25681 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n25682 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n25683 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n25684 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n25685 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n25686 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n25687 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n25688 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n25689 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n25690 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n25691 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n25692 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n25693 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n25694 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n25695 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n25696 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n25697 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n25698 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n25699 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n25700 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n25701 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n25702 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_1_3 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n25763 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n25764 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n25765 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n25766 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n25767 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n25768 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n25769 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n25770 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n25771 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n25772 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n25773 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n25774 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n25775 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n25776 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n25777 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n25778 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n25779 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n25780 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n25781 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n25782 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n25783 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n25829_o = {alu_7_i_n25602, alu_6_i_n25590, alu_5_i_n25578, alu_4_i_n25566, alu_3_i_n25554, alu_2_i_n25542, alu_1_i_n25530, alu_0_i_n25518};
  assign n25830_o = {alu_7_i_n25604, alu_6_i_n25592, alu_5_i_n25580, alu_4_i_n25568, alu_3_i_n25556, alu_2_i_n25544, alu_1_i_n25532, alu_0_i_n25520};
  assign n25831_o = {alu_7_i_n25603, alu_6_i_n25591, alu_5_i_n25579, alu_4_i_n25567, alu_3_i_n25555, alu_2_i_n25543, alu_1_i_n25531, alu_0_i_n25519};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25832_o = dp_readena_vm ? n25395_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25833_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n25833_q <= n25832_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25834_o = dp_readena_vm ? n25396_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25835_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n25835_q <= n25834_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25836_q <= 1'b0;
    else
      n25836_q <= n25407_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25837_q <= 1'b0;
    else
      n25837_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25838_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25839_q <= 1'b0;
    else
      n25839_q <= n25838_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25840_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25841_q <= 2'b00;
    else
      n25841_q <= n25840_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25842_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25843_q <= 2'b00;
    else
      n25843_q <= n25842_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25844_o = dp_readena_vm ? n25400_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25845_q <= 3'b000;
    else
      n25845_q <= n25844_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25846_o = dp_readena_vm ? n25402_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25847_q <= 3'b000;
    else
      n25847_q <= n25846_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25848_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25849_q <= 1'b0;
    else
      n25849_q <= n25848_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n25850_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n25343_o)
    if (n25343_o)
      n25851_q <= 2'b00;
    else
      n25851_q <= n25850_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25852_q <= 3'b000;
    else
      n25852_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25853_q <= 3'b000;
    else
      n25853_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25854_q <= 2'b00;
    else
      n25854_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25857_q <= 3'b000;
    else
      n25857_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25858_q <= 3'b000;
    else
      n25858_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25859_q <= 1'b0;
    else
      n25859_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25860_q <= 2'b00;
    else
      n25860_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25861_q <= 2'b00;
    else
      n25861_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25862_q <= 1'b0;
    else
      n25862_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25863_q <= 2'b00;
    else
      n25863_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25864_q <= 22'b0000000000000000000000;
    else
      n25864_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25865_q <= 3'b000;
    else
      n25865_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25866_q <= 22'b0000000000000000000000;
    else
      n25866_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25867_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n25867_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25868_o = n25016_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25869_q <= 1'b0;
    else
      n25869_q <= n25868_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25870_o = n25016_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25871_q <= 1'b0;
    else
      n25871_q <= n25870_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25872_o = n25162_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25873_q <= 1'b0;
    else
      n25873_q <= n25872_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25874_o = n25162_o ? dp_wr_fork : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25875_q <= 1'b0;
    else
      n25875_q <= n25874_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25876_q <= 22'b0000000000000000000000;
    else
      n25876_q <= n25014_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25877_q <= 22'b0000000000000000000000;
    else
      n25877_q <= n25160_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25878_o = n25162_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25879_q <= 6'b000000;
    else
      n25879_q <= n25878_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25880_o = n25162_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25881_q <= 1'b0;
    else
      n25881_q <= n25880_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25884_o = n25162_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25885_q <= 3'b000;
    else
      n25885_q <= n25884_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25886_o = n25162_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25887_q <= 2'b00;
    else
      n25887_q <= n25886_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25888_o = n25162_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25889_q <= 1'b0;
    else
      n25889_q <= n25888_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n25890_o = n25162_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25891_q <= 22'b0000000000000000000000;
    else
      n25891_q <= n25890_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25892_o = n25016_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25893_q <= 1'b0;
    else
      n25893_q <= n25892_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25894_o = n25016_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25895_q <= 3'b000;
    else
      n25895_q <= n25894_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25896_o = n25016_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25897_q <= 2'b00;
    else
      n25897_q <= n25896_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n25898_o = ~n25003_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n25899_o = n25016_o & n25898_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25900_o = n25899_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n25901_q <= n25900_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n25902_o = ~n25003_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n25903_o = n25016_o & n25902_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25904_o = n25903_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n25905_q <= n25904_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25906_o = n25016_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25907_q <= 1'b0;
    else
      n25907_q <= n25906_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25908_o = n25016_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25909_q <= 2'b00;
    else
      n25909_q <= n25908_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25910_o = n25016_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25911_q <= 2'b00;
    else
      n25911_q <= n25910_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25912_o = n25016_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25913_q <= 1'b0;
    else
      n25913_q <= n25912_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n25914_o = n25016_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25915_q <= 2'b00;
    else
      n25915_q <= n25914_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25916_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n25916_q <= n25174_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n25917_o = {n25217_o, n25916_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25918_q <= 3'b000;
    else
      n25918_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n25003_o)
    if (n25003_o)
      n25919_q <= 3'b000;
    else
      n25919_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n25149_o)
    if (n25149_o)
      n25920_q <= 3'b000;
    else
      n25920_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25922_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n25922_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25923_q <= 32'b00000000000000000000000000000000;
    else
      n25923_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25924_q <= 1'b0;
    else
      n25924_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25925_q <= 1'b0;
    else
      n25925_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25926_q <= 1'b0;
    else
      n25926_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25927_q <= 2'b00;
    else
      n25927_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25928_q <= 4'b0000;
    else
      n25928_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25929_q <= 1'b0;
    else
      n25929_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25930_q <= 4'b0000;
    else
      n25930_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25931_q <= 1'b0;
    else
      n25931_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25932_q <= 4'b0000;
    else
      n25932_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25933_q <= 1'b0;
    else
      n25933_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25934_q <= 1'b0;
    else
      n25934_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25935_q <= 2'b00;
    else
      n25935_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n25292_o)
    if (n25292_o)
      n25936_q <= 28'b0000000000000000000000000000;
    else
      n25936_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25937_q <= 1'b0;
    else
      n25937_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25938_q <= 1'b0;
    else
      n25938_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25940_q <= 1'b0;
    else
      n25940_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n25080_o)
    if (n25080_o)
      n25941_q <= 1'b0;
    else
      n25941_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25943_q <= 1'b0;
    else
      n25943_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25944_q <= 1'b0;
    else
      n25944_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25945_q <= 1'b0;
    else
      n25945_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25946_q <= 22'b0000000000000000000000;
    else
      n25946_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25947_q <= 1'b0;
    else
      n25947_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25948_q <= 22'b0000000000000000000000;
    else
      n25948_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25949_q <= 22'b0000000000000000000000;
    else
      n25949_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25950_q <= 1'b0;
    else
      n25950_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25951_q <= 22'b0000000000000000000000;
    else
      n25951_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25952_q <= 6'b000000;
    else
      n25952_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25953_q <= 1'b0;
    else
      n25953_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25954_q <= 1'b0;
    else
      n25954_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25955_q <= 1'b0;
    else
      n25955_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25956_q <= 3'b000;
    else
      n25956_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25957_q <= 2'b00;
    else
      n25957_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25958_q <= 1'b0;
    else
      n25958_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25959_q <= 1'b0;
    else
      n25959_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25960_q <= 3'b000;
    else
      n25960_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25961_q <= 2'b00;
    else
      n25961_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25962_q <= 1'b0;
    else
      n25962_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25963_q <= 2'b00;
    else
      n25963_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25964_q <= 2'b00;
    else
      n25964_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25965_q <= 1'b0;
    else
      n25965_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25966_q <= 2'b00;
    else
      n25966_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25967_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n25967_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n24807_o)
    if (n24807_o)
      n25968_q <= 1'b0;
    else
      n25968_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n25969_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n25970_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_1_2
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire dp_wr_fork;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire dp_wr_fork_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n23621_o;
  wire n23622_o;
  wire n23623_o;
  wire n23626_o;
  wire [4:0] n23714_o;
  wire n23715_o;
  wire [4:0] n23716_o;
  wire n23717_o;
  wire [2:0] n23720_o;
  wire [4:0] n23722_o;
  wire n23723_o;
  wire n23724_o;
  wire n23725_o;
  wire n23726_o;
  wire [4:0] n23727_o;
  wire [4:0] n23728_o;
  wire [4:0] n23729_o;
  wire n23730_o;
  wire n23731_o;
  wire n23732_o;
  wire [4:0] n23733_o;
  wire n23734_o;
  wire n23735_o;
  wire [4:0] n23736_o;
  wire n23737_o;
  wire n23738_o;
  wire n23739_o;
  wire n23740_o;
  wire n23743_o;
  wire n23749_o;
  wire n23751_o;
  wire [2:0] n23753_o;
  wire n23755_o;
  wire n23756_o;
  wire n23757_o;
  wire [2:0] n23759_o;
  wire [2:0] n23761_o;
  wire [2:0] n23763_o;
  wire n23764_o;
  wire n23765_o;
  wire [21:0] n23766_o;
  wire n23767_o;
  wire [2:0] n23768_o;
  wire [1:0] n23769_o;
  wire n23770_o;
  wire [21:0] n23771_o;
  wire n23772_o;
  wire [1:0] n23773_o;
  wire [1:0] n23774_o;
  wire n23775_o;
  wire [1:0] n23776_o;
  wire [2:0] n23777_o;
  wire [2:0] n23778_o;
  wire n23783_o;
  wire n23784_o;
  wire n23785_o;
  wire n23786_o;
  wire n23787_o;
  wire n23789_o;
  wire [2:0] n23791_o;
  wire n23793_o;
  wire n23794_o;
  wire n23795_o;
  wire [2:0] n23797_o;
  wire [2:0] n23801_o;
  wire [2:0] n23803_o;
  wire n23804_o;
  wire n23805_o;
  wire [21:0] n23806_o;
  wire [5:0] n23807_o;
  wire n23808_o;
  wire [2:0] n23809_o;
  wire [1:0] n23810_o;
  wire n23811_o;
  wire [21:0] n23812_o;
  wire [2:0] n23814_o;
  wire [2:0] n23817_o;
  wire n23822_o;
  wire n23825_o;
  wire n23826_o;
  wire [21:0] n23827_o;
  wire [21:0] n23829_o;
  wire [21:0] n23830_o;
  wire [21:0] n23832_o;
  wire [21:0] n23833_o;
  wire n23835_o;
  wire n23899_o;
  wire n23968_o;
  wire n23971_o;
  wire n23972_o;
  wire [21:0] n23973_o;
  wire [21:0] n23975_o;
  wire [21:0] n23976_o;
  wire [21:0] n23978_o;
  wire [21:0] n23979_o;
  wire n23981_o;
  wire [83:0] n23982_o;
  wire [83:0] n23983_o;
  wire [83:0] n23993_o;
  wire [11:0] n24035_o;
  wire [11:0] n24036_o;
  wire n24050_o;
  wire n24052_o;
  wire [11:0] n24053_o;
  wire [11:0] n24054_o;
  wire [11:0] n24055_o;
  wire [95:0] n24057_o;
  wire [95:0] n24058_o;
  wire [1:0] n24064_o;
  wire [2:0] n24065_o;
  wire n24066_o;
  wire n24068_o;
  wire n24069_o;
  wire n24071_o;
  wire n24072_o;
  wire n24075_o;
  wire n24077_o;
  wire n24078_o;
  wire n24081_o;
  wire n24082_o;
  wire [1:0] n24084_o;
  wire [1:0] n24086_o;
  wire n24088_o;
  wire [1:0] n24090_o;
  wire [1:0] n24096_o;
  wire [2:0] n24097_o;
  wire [4:0] n24098_o;
  wire n24101_o;
  wire [95:0] n24102_o;
  wire [95:0] n24104_o;
  wire n24106_o;
  wire n24111_o;
  wire n24162_o;
  wire n24165_o;
  wire [2:0] n24166_o;
  wire [11:0] n24167_o;
  wire n24169_o;
  wire [11:0] n24170_o;
  wire n24172_o;
  wire [11:0] n24173_o;
  wire n24175_o;
  wire [11:0] n24176_o;
  wire n24178_o;
  wire [11:0] n24179_o;
  wire n24181_o;
  wire [11:0] n24182_o;
  wire n24184_o;
  wire [11:0] n24185_o;
  wire n24187_o;
  wire [11:0] n24188_o;
  wire [6:0] n24189_o;
  wire [11:0] n24190_o;
  reg [11:0] n24191_o;
  wire [11:0] n24192_o;
  reg [11:0] n24193_o;
  wire [11:0] n24194_o;
  reg [11:0] n24195_o;
  wire [11:0] n24196_o;
  reg [11:0] n24197_o;
  wire [11:0] n24198_o;
  reg [11:0] n24199_o;
  wire [11:0] n24200_o;
  reg [11:0] n24201_o;
  wire [11:0] n24202_o;
  reg [11:0] n24203_o;
  wire [11:0] n24204_o;
  reg [11:0] n24205_o;
  wire n24207_o;
  wire n24210_o;
  wire [95:0] n24211_o;
  wire [95:0] n24212_o;
  wire [95:0] n24213_o;
  wire [95:0] n24214_o;
  wire [95:0] n24215_o;
  wire n24217_o;
  wire [2:0] n24219_o;
  wire [2:0] n24221_o;
  wire n24226_o;
  wire [12:0] xregister_file_i_n24275;
  wire [255:0] xregister_file_i_n24276;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n24281;
  wire [12:0] iregister_i_n24282;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n24289_o;
  wire n24291_o;
  wire n24292_o;
  wire n24294_o;
  wire n24295_o;
  wire n24298_o;
  wire n24300_o;
  wire n24301_o;
  wire n24304_o;
  wire n24305_o;
  wire [4:0] n24313_o;
  wire n24314_o;
  wire [4:0] n24315_o;
  wire [4:0] n24318_o;
  wire [4:0] n24319_o;
  wire [4:0] n24320_o;
  wire n24321_o;
  wire n24322_o;
  wire n24323_o;
  wire n24324_o;
  wire n24325_o;
  wire n24326_o;
  wire n24327_o;
  wire n24328_o;
  wire n24329_o;
  wire n24332_o;
  wire [31:0] n24334_o;
  wire [11:0] n24335_o;
  wire [11:0] n24336_o;
  wire [31:0] alu_0_i_n24337;
  wire alu_0_i_n24338;
  wire [11:0] alu_0_i_n24339;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n24346_o;
  wire [11:0] n24347_o;
  wire [11:0] n24348_o;
  wire [31:0] alu_1_i_n24349;
  wire alu_1_i_n24350;
  wire [11:0] alu_1_i_n24351;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n24358_o;
  wire [11:0] n24359_o;
  wire [11:0] n24360_o;
  wire [31:0] alu_2_i_n24361;
  wire alu_2_i_n24362;
  wire [11:0] alu_2_i_n24363;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n24370_o;
  wire [11:0] n24371_o;
  wire [11:0] n24372_o;
  wire [31:0] alu_3_i_n24373;
  wire alu_3_i_n24374;
  wire [11:0] alu_3_i_n24375;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n24382_o;
  wire [11:0] n24383_o;
  wire [11:0] n24384_o;
  wire [31:0] alu_4_i_n24385;
  wire alu_4_i_n24386;
  wire [11:0] alu_4_i_n24387;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n24394_o;
  wire [11:0] n24395_o;
  wire [11:0] n24396_o;
  wire [31:0] alu_5_i_n24397;
  wire alu_5_i_n24398;
  wire [11:0] alu_5_i_n24399;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n24406_o;
  wire [11:0] n24407_o;
  wire [11:0] n24408_o;
  wire [31:0] alu_6_i_n24409;
  wire alu_6_i_n24410;
  wire [11:0] alu_6_i_n24411;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n24418_o;
  wire [11:0] n24419_o;
  wire [11:0] n24420_o;
  wire [31:0] alu_7_i_n24421;
  wire alu_7_i_n24422;
  wire [11:0] alu_7_i_n24423;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n24430_o;
  wire n24431_o;
  wire [12:0] ialu_i_n24432;
  wire ialu_i_n24433;
  wire ialu_i_n24434;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n24443;
  wire [95:0] register_bank_i_n24444;
  wire [16:0] n24445_o;
  wire [16:0] n24446_o;
  wire [95:0] register_bank_i_n24447;
  wire register_bank_i_n24448;
  wire register_bank_i_n24449;
  wire [2:0] register_bank_i_n24450;
  wire [2:0] register_bank_i_n24451;
  wire [1:0] register_bank_i_n24452;
  wire [2:0] register_bank_i_n24453;
  wire [2:0] register_bank_i_n24454;
  wire register_bank_i_n24455;
  wire [1:0] register_bank_i_n24456;
  wire [1:0] register_bank_i_n24457;
  wire register_bank_i_n24458;
  wire [1:0] register_bank_i_n24459;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n24492;
  wire instr_decoder2_i_n24493;
  wire [3:0] instr_decoder2_i_n24494;
  wire instr_decoder2_i_n24495;
  wire instr_decoder2_i_n24496;
  wire instr_decoder2_i_n24497;
  wire instr_decoder2_i_n24498;
  wire [11:0] instr_decoder2_i_n24499;
  wire [11:0] instr_decoder2_i_n24500;
  wire [11:0] instr_decoder2_i_n24501;
  wire instr_decoder2_i_n24502;
  wire instr_decoder2_i_n24503;
  wire instr_decoder2_i_n24504;
  wire [7:0] instr_decoder2_i_n24505;
  wire instr_decoder2_i_n24506;
  wire [11:0] instr_decoder2_i_n24507;
  wire instr_decoder2_i_n24508;
  wire instr_decoder2_i_n24509;
  wire [3:0] instr_decoder2_i_n24510;
  wire [3:0] instr_decoder2_i_n24511;
  wire instr_decoder2_i_n24512;
  wire instr_decoder2_i_n24513;
  wire [2:0] instr_decoder2_i_n24514;
  wire [12:0] instr_decoder2_i_n24515;
  wire instr_decoder2_i_n24516;
  wire [4:0] instr_decoder2_i_n24517;
  wire [12:0] instr_decoder2_i_n24518;
  wire [12:0] instr_decoder2_i_n24519;
  wire [7:0] instr_decoder2_i_n24520;
  wire [7:0] instr_decoder2_i_n24521;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n24582;
  wire instr_dispatch2_i1_n24583;
  wire [11:0] instr_dispatch2_i1_n24584;
  wire [11:0] instr_dispatch2_i1_n24585;
  wire instr_dispatch2_i1_n24586;
  wire instr_dispatch2_i1_n24587;
  wire instr_dispatch2_i1_n24588;
  wire instr_dispatch2_i1_n24589;
  wire instr_dispatch2_i1_n24590;
  wire instr_dispatch2_i1_n24591;
  wire instr_dispatch2_i1_n24592;
  wire instr_dispatch2_i1_n24593;
  wire [11:0] instr_dispatch2_i1_n24594;
  wire [7:0] instr_dispatch2_i1_n24595;
  wire [95:0] instr_dispatch2_i1_n24596;
  wire [7:0] instr_dispatch2_i1_n24597;
  wire [95:0] instr_dispatch2_i1_n24598;
  wire [95:0] instr_dispatch2_i1_n24599;
  wire [11:0] instr_dispatch2_i1_n24600;
  wire [4:0] instr_dispatch2_i1_n24601;
  wire [3:0] instr_dispatch2_i1_n24602;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n24648_o;
  wire [95:0] n24649_o;
  wire [7:0] n24650_o;
  wire [95:0] n24651_o;
  reg [95:0] n24652_q;
  wire [95:0] n24653_o;
  reg [95:0] n24654_q;
  reg n24655_q;
  reg n24656_q;
  wire n24657_o;
  reg n24658_q;
  wire [1:0] n24659_o;
  reg [1:0] n24660_q;
  wire [1:0] n24661_o;
  reg [1:0] n24662_q;
  wire [2:0] n24663_o;
  reg [2:0] n24664_q;
  wire [2:0] n24665_o;
  reg [2:0] n24666_q;
  wire n24667_o;
  reg n24668_q;
  wire [1:0] n24669_o;
  reg [1:0] n24670_q;
  reg [2:0] n24671_q;
  reg [2:0] n24672_q;
  reg [1:0] n24673_q;
  reg [2:0] n24676_q;
  reg [2:0] n24677_q;
  reg n24678_q;
  reg [1:0] n24679_q;
  reg [1:0] n24680_q;
  reg n24681_q;
  reg [1:0] n24682_q;
  reg [21:0] n24683_q;
  reg [2:0] n24684_q;
  reg [21:0] n24685_q;
  reg [95:0] n24686_q;
  wire n24687_o;
  reg n24688_q;
  wire n24689_o;
  reg n24690_q;
  wire n24691_o;
  reg n24692_q;
  wire n24693_o;
  reg n24694_q;
  reg [21:0] n24695_q;
  reg [21:0] n24696_q;
  wire [5:0] n24697_o;
  reg [5:0] n24698_q;
  wire n24699_o;
  reg n24700_q;
  wire [2:0] n24703_o;
  reg [2:0] n24704_q;
  wire [1:0] n24705_o;
  reg [1:0] n24706_q;
  wire n24707_o;
  reg n24708_q;
  wire [21:0] n24709_o;
  reg [21:0] n24710_q;
  wire n24711_o;
  reg n24712_q;
  wire [2:0] n24713_o;
  reg [2:0] n24714_q;
  wire [1:0] n24715_o;
  reg [1:0] n24716_q;
  wire n24717_o;
  wire n24718_o;
  wire n24719_o;
  reg n24720_q;
  wire n24721_o;
  wire n24722_o;
  wire [21:0] n24723_o;
  reg [21:0] n24724_q;
  wire n24725_o;
  reg n24726_q;
  wire [1:0] n24727_o;
  reg [1:0] n24728_q;
  wire [1:0] n24729_o;
  reg [1:0] n24730_q;
  wire n24731_o;
  reg n24732_q;
  wire [1:0] n24733_o;
  reg [1:0] n24734_q;
  reg [83:0] n24735_q;
  wire [95:0] n24736_o;
  reg [2:0] n24737_q;
  reg [2:0] n24738_q;
  reg [2:0] n24739_q;
  reg [79:0] n24741_q;
  reg [31:0] n24742_q;
  reg n24743_q;
  reg n24744_q;
  reg n24745_q;
  reg [1:0] n24746_q;
  reg [3:0] n24747_q;
  reg n24748_q;
  reg [3:0] n24749_q;
  reg n24750_q;
  reg [3:0] n24751_q;
  reg n24752_q;
  reg n24753_q;
  reg [1:0] n24754_q;
  reg [27:0] n24755_q;
  reg n24756_q;
  reg n24757_q;
  reg n24759_q;
  reg n24760_q;
  reg n24762_q;
  reg n24763_q;
  reg n24764_q;
  reg [21:0] n24765_q;
  reg n24766_q;
  reg [21:0] n24767_q;
  reg [21:0] n24768_q;
  reg n24769_q;
  reg [21:0] n24770_q;
  reg [5:0] n24771_q;
  reg n24772_q;
  reg n24773_q;
  reg n24774_q;
  reg [2:0] n24775_q;
  reg [1:0] n24776_q;
  reg n24777_q;
  reg n24778_q;
  reg [2:0] n24779_q;
  reg [1:0] n24780_q;
  reg n24781_q;
  reg [1:0] n24782_q;
  reg [1:0] n24783_q;
  reg n24784_q;
  reg [1:0] n24785_q;
  reg [95:0] n24786_q;
  reg n24787_q;
  wire [2:0] n24788_o;
  wire [2:0] n24789_o;
  assign i_y_neg_out = n24430_o;
  assign i_y_zero_out = n24431_o;
  assign dp_readdata_out = n24104_o;
  assign dp_readdata_vm_out = n24106_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n24788_o;
  assign dp_read_vaddr_out = n24789_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n24084_o;
  assign dp_read_data_type_out = n24086_o;
  assign dp_read_stream_out = n24088_o;
  assign dp_read_stream_id_out = n24090_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n24443; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n24444; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n24582; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n24583; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n24591; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n24588; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n24589; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n24590; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n24596; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n24597; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n24499; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n24500; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n24501; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n24282; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n24516; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n24492; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n24598; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n24599; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n24600; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n24648_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n24649_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n24650_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n24601; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n24602; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n24494; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n24332_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n24305_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n24098_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n24584; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n24585; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n24594; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n24595; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n24096_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n24097_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n24493; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n24498; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n24495; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n24496; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n24497; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n24506; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n24507; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n24502; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n24503; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n24504; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n24505; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n24586; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n24587; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n24593; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n24508; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n24509; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n24510; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n24281; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n24511; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n24512; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n24513; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n24514; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n24515; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n24652_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n24654_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n24655_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n24656_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n24658_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n24660_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n24662_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n24664_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n24666_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n24668_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n24670_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n24517; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n24518; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n24519; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n24432; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n24433; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n24434; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n24592; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n24520; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n24521; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n24275; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n24276; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n23764_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n23765_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n23804_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:191:8  */
  assign dp_wr_fork = n23805_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n23766_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n23806_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n23807_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n23808_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n23809_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n23810_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n23811_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n23812_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n23767_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n23768_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n23769_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n23770_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n23771_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n23772_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n23773_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n23774_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n23775_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n23776_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n24058_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n23777_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n23778_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n23814_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n23817_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n24671_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n24672_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n24673_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n24676_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n24677_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n24678_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n24679_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n24680_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n24681_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n24682_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n24683_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n24684_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n24685_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n24686_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n24688_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n24690_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n24692_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:238:8  */
  assign dp_wr_fork_r = n24694_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n24695_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n24696_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n24698_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n24700_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n24704_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n24706_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n24708_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n24710_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n24712_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n24714_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n24716_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n24720_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n24724_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n24726_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n24728_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n24730_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n24732_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n24734_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n24736_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n24737_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n24738_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n24739_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n24082_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n23743_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n24449; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n24450; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n24451; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n24452; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n24453; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n24454; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n24447; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n24448; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n24455; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n24456; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n24457; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n24458; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n24459; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n23621_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n23622_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n23623_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n24741_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n24742_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n24743_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n24744_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n24745_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n24746_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n24747_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n24748_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n24749_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n24750_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n24751_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n24752_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n24753_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n24754_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n24755_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n24756_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n24757_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n24759_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n24760_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n24762_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n24763_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n24764_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n24765_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n24766_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n24767_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n24768_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n24769_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n24770_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n24771_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n24772_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n24773_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n24774_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n24775_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n24776_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n24777_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n24778_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n24779_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n24780_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n24781_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n24782_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n24783_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n24784_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n24785_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n24786_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n24787_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n23621_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n23622_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n23623_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n23626_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n23714_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n23715_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n23716_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n23717_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n23720_o = n23717_o ? 3'b001 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n23722_o = n23716_o + n23714_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n23723_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n23724_o = n23723_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n23725_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n23726_o = n23725_o & n23724_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n23727_o = n23714_o & n23716_o;
  /* ../../HW/src/pcore/pcore.vhd:104:8  */
  assign n23728_o = {n23720_o, 2'b10};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n23729_o = n23714_o & n23728_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n23730_o = n23727_o == n23729_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n23731_o = n23730_o & n23715_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n23732_o = ~n23715_o;
  /* ../../HW/src/pcore/pcore.vhd:349:1  */
  assign n23733_o = {n23720_o, 2'b10};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n23734_o = $unsigned(n23733_o) >= $unsigned(n23716_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n23735_o = n23734_o & n23732_o;
  /* ../../HW/src/pcore/pcore.vhd:349:1  */
  assign n23736_o = {n23720_o, 2'b10};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n23737_o = $unsigned(n23736_o) <= $unsigned(n23722_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n23738_o = n23737_o & n23735_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n23739_o = n23731_o | n23738_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n23740_o = n23739_o & n23726_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n23743_o = n23740_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n23749_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n23751_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n23753_o = n23751_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n23755_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n23756_o = n23755_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n23757_o = dp_read_gen_valid_in_r & n23756_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n23759_o = n23757_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n23761_o = n23757_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n23763_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23764_o = n23749_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23765_o = n23749_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23766_o = n23749_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23767_o = n23749_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23768_o = n23749_o ? n23753_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23769_o = n23749_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23770_o = n23749_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23771_o = n23749_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23772_o = n23749_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23773_o = n23749_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23774_o = n23749_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23775_o = n23749_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23776_o = n23749_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23777_o = n23749_o ? n23759_o : n23763_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n23778_o = n23749_o ? n23761_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n23783_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n23784_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n23785_o = dp_write_in_r & n23784_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n23786_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n23787_o = n23785_o & n23786_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n23789_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n23791_o = n23789_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n23793_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n23794_o = n23793_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n23795_o = dp_write_gen_valid_in_r & n23794_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n23797_o = n23795_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n23801_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n23803_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23804_o = n23783_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23805_o = n23783_o ? dp_wr_fork_in_r : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23806_o = n23783_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23807_o = n23783_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23808_o = n23783_o ? n23787_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23809_o = n23783_o ? n23791_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23810_o = n23783_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23811_o = n23783_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23812_o = n23783_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23814_o = n23783_o ? n23797_o : n23801_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n23817_o = n23783_o ? 3'b000 : n23803_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n23822_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n23825_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n23826_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n23827_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n23829_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n23830_o = n23826_o ? n23827_o : n23829_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n23832_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n23833_o = n23825_o ? n23830_o : n23832_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n23835_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n23899_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n23968_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n23971_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n23972_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n23973_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n23975_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n23976_o = n23972_o ? n23973_o : n23975_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n23978_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n23979_o = n23971_o ? n23976_o : n23978_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n23981_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n23982_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n23983_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n23993_o = n23981_o ? n23982_o : n23983_o;
  assign n24035_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n24036_o = n23968_o ? 12'b000000000000 : n24035_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n24050_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n24052_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n24053_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n24054_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n24055_o = n24052_o ? n24053_o : n24054_o;
  assign n24057_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n24055_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n24058_o = n24050_o ? n24057_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n24064_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n24065_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n24066_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n24068_o = n24064_o == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n24069_o = n24068_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n24071_o = n24065_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n24072_o = n24071_o & n24069_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n24075_o = n24072_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n24077_o = n24064_o == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n24078_o = n24077_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n24081_o = n24078_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n24082_o = n24066_o ? n24075_o : n24081_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n24084_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n24086_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n24088_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n24090_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n24096_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n24097_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n24098_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n24101_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n24102_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n24104_o = n24101_o ? 96'bZ : n24102_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n24106_o = n24101_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n24111_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n24162_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n24165_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n24166_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n24167_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n24169_o = n24166_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n24170_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n24172_o = n24166_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n24173_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n24175_o = n24166_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n24176_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n24178_o = n24166_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n24179_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n24181_o = n24166_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n24182_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n24184_o = n24166_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n24185_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n24187_o = n24166_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n24188_o = dp_readdata_vm[11:0];
  assign n24189_o = {n24187_o, n24184_o, n24181_o, n24178_o, n24175_o, n24172_o, n24169_o};
  assign n24190_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24191_o = n24190_o;
      7'b0100000: n24191_o = n24190_o;
      7'b0010000: n24191_o = n24190_o;
      7'b0001000: n24191_o = n24190_o;
      7'b0000100: n24191_o = n24190_o;
      7'b0000010: n24191_o = n24190_o;
      7'b0000001: n24191_o = n24190_o;
      default: n24191_o = n24188_o;
    endcase
  assign n24192_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24193_o = n24185_o;
      7'b0100000: n24193_o = n24192_o;
      7'b0010000: n24193_o = n24192_o;
      7'b0001000: n24193_o = n24192_o;
      7'b0000100: n24193_o = n24192_o;
      7'b0000010: n24193_o = n24192_o;
      7'b0000001: n24193_o = n24192_o;
      default: n24193_o = n24192_o;
    endcase
  assign n24194_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24195_o = n24194_o;
      7'b0100000: n24195_o = n24182_o;
      7'b0010000: n24195_o = n24194_o;
      7'b0001000: n24195_o = n24194_o;
      7'b0000100: n24195_o = n24194_o;
      7'b0000010: n24195_o = n24194_o;
      7'b0000001: n24195_o = n24194_o;
      default: n24195_o = n24194_o;
    endcase
  assign n24196_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24197_o = n24196_o;
      7'b0100000: n24197_o = n24196_o;
      7'b0010000: n24197_o = n24179_o;
      7'b0001000: n24197_o = n24196_o;
      7'b0000100: n24197_o = n24196_o;
      7'b0000010: n24197_o = n24196_o;
      7'b0000001: n24197_o = n24196_o;
      default: n24197_o = n24196_o;
    endcase
  assign n24198_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24199_o = n24198_o;
      7'b0100000: n24199_o = n24198_o;
      7'b0010000: n24199_o = n24198_o;
      7'b0001000: n24199_o = n24176_o;
      7'b0000100: n24199_o = n24198_o;
      7'b0000010: n24199_o = n24198_o;
      7'b0000001: n24199_o = n24198_o;
      default: n24199_o = n24198_o;
    endcase
  assign n24200_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24201_o = n24200_o;
      7'b0100000: n24201_o = n24200_o;
      7'b0010000: n24201_o = n24200_o;
      7'b0001000: n24201_o = n24200_o;
      7'b0000100: n24201_o = n24173_o;
      7'b0000010: n24201_o = n24200_o;
      7'b0000001: n24201_o = n24200_o;
      default: n24201_o = n24200_o;
    endcase
  assign n24202_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24203_o = n24202_o;
      7'b0100000: n24203_o = n24202_o;
      7'b0010000: n24203_o = n24202_o;
      7'b0001000: n24203_o = n24202_o;
      7'b0000100: n24203_o = n24202_o;
      7'b0000010: n24203_o = n24170_o;
      7'b0000001: n24203_o = n24202_o;
      default: n24203_o = n24202_o;
    endcase
  assign n24204_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n24189_o)
      7'b1000000: n24205_o = n24204_o;
      7'b0100000: n24205_o = n24204_o;
      7'b0010000: n24205_o = n24204_o;
      7'b0001000: n24205_o = n24204_o;
      7'b0000100: n24205_o = n24204_o;
      7'b0000010: n24205_o = n24204_o;
      7'b0000001: n24205_o = n24167_o;
      default: n24205_o = n24204_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n24207_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n24210_o = n24207_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n24211_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n24212_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n24213_o = {n24205_o, n24203_o, n24201_o, n24199_o, n24197_o, n24195_o, n24193_o, n24191_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n24214_o = n24165_o ? n24213_o : n24211_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n24215_o = n24165_o ? dp_readdata2_r : n24212_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n24217_o = n24165_o ? n24210_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n24219_o = n24165_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n24221_o = n24165_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n24226_o = dp_readena_vm ? n24217_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n24275 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n24276 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n24281 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n24282 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n24289_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n24291_o = dp_rd_pid == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n24292_o = n24291_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n24294_o = dp_rd_cid == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n24295_o = n24294_o & n24292_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n24298_o = n24295_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n24300_o = dp_rd_pid == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n24301_o = n24300_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n24304_o = n24301_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n24305_o = n24289_o ? n24298_o : n24304_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n24313_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n24314_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n24315_o = dp_mcast_addr + n24313_o;
  /* ../../HW/src/pcore/pcore.vhd:1022:1  */
  assign n24318_o = dp_wr_fork ? 5'b00010 : 5'b00110;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n24319_o = n24313_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n24320_o = n24313_o & n24318_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n24321_o = n24319_o == n24320_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n24322_o = n24321_o & n24314_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n24323_o = ~n24314_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n24324_o = $unsigned(n24318_o) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n24325_o = n24324_o & n24323_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n24326_o = $unsigned(n24318_o) <= $unsigned(n24315_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n24327_o = n24326_o & n24325_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n24328_o = n24322_o | n24327_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n24329_o = n24328_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n24332_o = n24329_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n24334_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n24335_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n24336_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n24337 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n24338 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n24339 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24334_o),
    .x1_in(n24335_o),
    .x2_in(n24336_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n24346_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n24347_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n24348_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n24349 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n24350 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n24351 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24346_o),
    .x1_in(n24347_o),
    .x2_in(n24348_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n24358_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n24359_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n24360_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n24361 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n24362 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n24363 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24358_o),
    .x1_in(n24359_o),
    .x2_in(n24360_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n24370_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n24371_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n24372_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n24373 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n24374 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n24375 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24370_o),
    .x1_in(n24371_o),
    .x2_in(n24372_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n24382_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n24383_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n24384_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n24385 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n24386 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n24387 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24382_o),
    .x1_in(n24383_o),
    .x2_in(n24384_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n24394_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n24395_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n24396_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n24397 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n24398 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n24399 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24394_o),
    .x1_in(n24395_o),
    .x2_in(n24396_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n24406_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n24407_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n24408_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n24409 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n24410 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n24411 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24406_o),
    .x1_in(n24407_o),
    .x2_in(n24408_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n24418_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n24419_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n24420_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n24421 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n24422 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n24423 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n24418_o),
    .x1_in(n24419_o),
    .x2_in(n24420_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n24430_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n24431_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n24432 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n24433 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n24434 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n24443 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n24444 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n24445_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n24446_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n24447 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n24448 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n24449 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n24450 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n24451 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n24452 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n24453 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n24454 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n24455 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n24456 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n24457 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n24458 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n24459 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n24445_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n24446_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n24492 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n24493 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n24494 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n24495 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n24496 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n24497 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n24498 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n24499 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n24500 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n24501 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n24502 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n24503 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n24504 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n24505 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n24506 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n24507 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n24508 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n24509 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n24510 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n24511 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n24512 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n24513 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n24514 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n24515 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n24516 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n24517 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n24518 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n24519 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n24520 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n24521 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_1_2 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n24582 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n24583 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n24584 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n24585 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n24586 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n24587 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n24588 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n24589 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n24590 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n24591 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n24592 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n24593 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n24594 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n24595 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n24596 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n24597 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n24598 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n24599 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n24600 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n24601 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n24602 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n24648_o = {alu_7_i_n24421, alu_6_i_n24409, alu_5_i_n24397, alu_4_i_n24385, alu_3_i_n24373, alu_2_i_n24361, alu_1_i_n24349, alu_0_i_n24337};
  assign n24649_o = {alu_7_i_n24423, alu_6_i_n24411, alu_5_i_n24399, alu_4_i_n24387, alu_3_i_n24375, alu_2_i_n24363, alu_1_i_n24351, alu_0_i_n24339};
  assign n24650_o = {alu_7_i_n24422, alu_6_i_n24410, alu_5_i_n24398, alu_4_i_n24386, alu_3_i_n24374, alu_2_i_n24362, alu_1_i_n24350, alu_0_i_n24338};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24651_o = dp_readena_vm ? n24214_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24652_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n24652_q <= n24651_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24653_o = dp_readena_vm ? n24215_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24654_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n24654_q <= n24653_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24655_q <= 1'b0;
    else
      n24655_q <= n24226_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24656_q <= 1'b0;
    else
      n24656_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24657_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24658_q <= 1'b0;
    else
      n24658_q <= n24657_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24659_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24660_q <= 2'b00;
    else
      n24660_q <= n24659_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24661_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24662_q <= 2'b00;
    else
      n24662_q <= n24661_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24663_o = dp_readena_vm ? n24219_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24664_q <= 3'b000;
    else
      n24664_q <= n24663_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24665_o = dp_readena_vm ? n24221_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24666_q <= 3'b000;
    else
      n24666_q <= n24665_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24667_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24668_q <= 1'b0;
    else
      n24668_q <= n24667_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n24669_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n24162_o)
    if (n24162_o)
      n24670_q <= 2'b00;
    else
      n24670_q <= n24669_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24671_q <= 3'b000;
    else
      n24671_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24672_q <= 3'b000;
    else
      n24672_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24673_q <= 2'b00;
    else
      n24673_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24676_q <= 3'b000;
    else
      n24676_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24677_q <= 3'b000;
    else
      n24677_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24678_q <= 1'b0;
    else
      n24678_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24679_q <= 2'b00;
    else
      n24679_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24680_q <= 2'b00;
    else
      n24680_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24681_q <= 1'b0;
    else
      n24681_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24682_q <= 2'b00;
    else
      n24682_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24683_q <= 22'b0000000000000000000000;
    else
      n24683_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24684_q <= 3'b000;
    else
      n24684_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24685_q <= 22'b0000000000000000000000;
    else
      n24685_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24686_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n24686_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24687_o = n23835_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24688_q <= 1'b0;
    else
      n24688_q <= n24687_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24689_o = n23835_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24690_q <= 1'b0;
    else
      n24690_q <= n24689_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24691_o = n23981_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24692_q <= 1'b0;
    else
      n24692_q <= n24691_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24693_o = n23981_o ? dp_wr_fork : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24694_q <= 1'b0;
    else
      n24694_q <= n24693_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24695_q <= 22'b0000000000000000000000;
    else
      n24695_q <= n23833_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24696_q <= 22'b0000000000000000000000;
    else
      n24696_q <= n23979_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24697_o = n23981_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24698_q <= 6'b000000;
    else
      n24698_q <= n24697_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24699_o = n23981_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24700_q <= 1'b0;
    else
      n24700_q <= n24699_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24703_o = n23981_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24704_q <= 3'b000;
    else
      n24704_q <= n24703_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24705_o = n23981_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24706_q <= 2'b00;
    else
      n24706_q <= n24705_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24707_o = n23981_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24708_q <= 1'b0;
    else
      n24708_q <= n24707_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n24709_o = n23981_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24710_q <= 22'b0000000000000000000000;
    else
      n24710_q <= n24709_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24711_o = n23835_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24712_q <= 1'b0;
    else
      n24712_q <= n24711_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24713_o = n23835_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24714_q <= 3'b000;
    else
      n24714_q <= n24713_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24715_o = n23835_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24716_q <= 2'b00;
    else
      n24716_q <= n24715_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n24717_o = ~n23822_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n24718_o = n23835_o & n24717_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24719_o = n24718_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n24720_q <= n24719_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n24721_o = ~n23822_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n24722_o = n23835_o & n24721_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24723_o = n24722_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n24724_q <= n24723_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24725_o = n23835_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24726_q <= 1'b0;
    else
      n24726_q <= n24725_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24727_o = n23835_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24728_q <= 2'b00;
    else
      n24728_q <= n24727_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24729_o = n23835_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24730_q <= 2'b00;
    else
      n24730_q <= n24729_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24731_o = n23835_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24732_q <= 1'b0;
    else
      n24732_q <= n24731_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n24733_o = n23835_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24734_q <= 2'b00;
    else
      n24734_q <= n24733_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24735_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n24735_q <= n23993_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n24736_o = {n24036_o, n24735_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24737_q <= 3'b000;
    else
      n24737_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n23822_o)
    if (n23822_o)
      n24738_q <= 3'b000;
    else
      n24738_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n23968_o)
    if (n23968_o)
      n24739_q <= 3'b000;
    else
      n24739_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24741_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n24741_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24742_q <= 32'b00000000000000000000000000000000;
    else
      n24742_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24743_q <= 1'b0;
    else
      n24743_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24744_q <= 1'b0;
    else
      n24744_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24745_q <= 1'b0;
    else
      n24745_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24746_q <= 2'b00;
    else
      n24746_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24747_q <= 4'b0000;
    else
      n24747_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24748_q <= 1'b0;
    else
      n24748_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24749_q <= 4'b0000;
    else
      n24749_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24750_q <= 1'b0;
    else
      n24750_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24751_q <= 4'b0000;
    else
      n24751_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24752_q <= 1'b0;
    else
      n24752_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24753_q <= 1'b0;
    else
      n24753_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24754_q <= 2'b00;
    else
      n24754_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n24111_o)
    if (n24111_o)
      n24755_q <= 28'b0000000000000000000000000000;
    else
      n24755_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24756_q <= 1'b0;
    else
      n24756_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24757_q <= 1'b0;
    else
      n24757_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24759_q <= 1'b0;
    else
      n24759_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n23899_o)
    if (n23899_o)
      n24760_q <= 1'b0;
    else
      n24760_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24762_q <= 1'b0;
    else
      n24762_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24763_q <= 1'b0;
    else
      n24763_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24764_q <= 1'b0;
    else
      n24764_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24765_q <= 22'b0000000000000000000000;
    else
      n24765_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24766_q <= 1'b0;
    else
      n24766_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24767_q <= 22'b0000000000000000000000;
    else
      n24767_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24768_q <= 22'b0000000000000000000000;
    else
      n24768_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24769_q <= 1'b0;
    else
      n24769_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24770_q <= 22'b0000000000000000000000;
    else
      n24770_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24771_q <= 6'b000000;
    else
      n24771_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24772_q <= 1'b0;
    else
      n24772_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24773_q <= 1'b0;
    else
      n24773_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24774_q <= 1'b0;
    else
      n24774_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24775_q <= 3'b000;
    else
      n24775_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24776_q <= 2'b00;
    else
      n24776_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24777_q <= 1'b0;
    else
      n24777_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24778_q <= 1'b0;
    else
      n24778_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24779_q <= 3'b000;
    else
      n24779_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24780_q <= 2'b00;
    else
      n24780_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24781_q <= 1'b0;
    else
      n24781_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24782_q <= 2'b00;
    else
      n24782_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24783_q <= 2'b00;
    else
      n24783_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24784_q <= 1'b0;
    else
      n24784_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24785_q <= 2'b00;
    else
      n24785_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24786_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n24786_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n23626_o)
    if (n23626_o)
      n24787_q <= 1'b0;
    else
      n24787_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n24788_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n24789_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_1_1
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire dp_wr_fork;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire dp_wr_fork_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n22440_o;
  wire n22441_o;
  wire n22442_o;
  wire n22445_o;
  wire [4:0] n22533_o;
  wire n22534_o;
  wire [4:0] n22535_o;
  wire n22536_o;
  wire [2:0] n22539_o;
  wire [4:0] n22541_o;
  wire n22542_o;
  wire n22543_o;
  wire n22544_o;
  wire n22545_o;
  wire [4:0] n22546_o;
  wire [4:0] n22547_o;
  wire [4:0] n22548_o;
  wire n22549_o;
  wire n22550_o;
  wire n22551_o;
  wire [4:0] n22552_o;
  wire n22553_o;
  wire n22554_o;
  wire [4:0] n22555_o;
  wire n22556_o;
  wire n22557_o;
  wire n22558_o;
  wire n22559_o;
  wire n22562_o;
  wire n22568_o;
  wire n22570_o;
  wire [2:0] n22572_o;
  wire n22574_o;
  wire n22575_o;
  wire n22576_o;
  wire [2:0] n22578_o;
  wire [2:0] n22580_o;
  wire [2:0] n22582_o;
  wire n22583_o;
  wire n22584_o;
  wire [21:0] n22585_o;
  wire n22586_o;
  wire [2:0] n22587_o;
  wire [1:0] n22588_o;
  wire n22589_o;
  wire [21:0] n22590_o;
  wire n22591_o;
  wire [1:0] n22592_o;
  wire [1:0] n22593_o;
  wire n22594_o;
  wire [1:0] n22595_o;
  wire [2:0] n22596_o;
  wire [2:0] n22597_o;
  wire n22602_o;
  wire n22603_o;
  wire n22604_o;
  wire n22605_o;
  wire n22606_o;
  wire n22608_o;
  wire [2:0] n22610_o;
  wire n22612_o;
  wire n22613_o;
  wire n22614_o;
  wire [2:0] n22616_o;
  wire [2:0] n22620_o;
  wire [2:0] n22622_o;
  wire n22623_o;
  wire n22624_o;
  wire [21:0] n22625_o;
  wire [5:0] n22626_o;
  wire n22627_o;
  wire [2:0] n22628_o;
  wire [1:0] n22629_o;
  wire n22630_o;
  wire [21:0] n22631_o;
  wire [2:0] n22633_o;
  wire [2:0] n22636_o;
  wire n22641_o;
  wire n22644_o;
  wire n22645_o;
  wire [21:0] n22646_o;
  wire [21:0] n22648_o;
  wire [21:0] n22649_o;
  wire [21:0] n22651_o;
  wire [21:0] n22652_o;
  wire n22654_o;
  wire n22718_o;
  wire n22787_o;
  wire n22790_o;
  wire n22791_o;
  wire [21:0] n22792_o;
  wire [21:0] n22794_o;
  wire [21:0] n22795_o;
  wire [21:0] n22797_o;
  wire [21:0] n22798_o;
  wire n22800_o;
  wire [83:0] n22801_o;
  wire [83:0] n22802_o;
  wire [83:0] n22812_o;
  wire [11:0] n22854_o;
  wire [11:0] n22855_o;
  wire n22869_o;
  wire n22871_o;
  wire [11:0] n22872_o;
  wire [11:0] n22873_o;
  wire [11:0] n22874_o;
  wire [95:0] n22876_o;
  wire [95:0] n22877_o;
  wire [1:0] n22883_o;
  wire [2:0] n22884_o;
  wire n22885_o;
  wire n22887_o;
  wire n22888_o;
  wire n22890_o;
  wire n22891_o;
  wire n22894_o;
  wire n22896_o;
  wire n22897_o;
  wire n22900_o;
  wire n22901_o;
  wire [1:0] n22903_o;
  wire [1:0] n22905_o;
  wire n22907_o;
  wire [1:0] n22909_o;
  wire [1:0] n22915_o;
  wire [2:0] n22916_o;
  wire [4:0] n22917_o;
  wire n22920_o;
  wire [95:0] n22921_o;
  wire [95:0] n22923_o;
  wire n22925_o;
  wire n22930_o;
  wire n22981_o;
  wire n22984_o;
  wire [2:0] n22985_o;
  wire [11:0] n22986_o;
  wire n22988_o;
  wire [11:0] n22989_o;
  wire n22991_o;
  wire [11:0] n22992_o;
  wire n22994_o;
  wire [11:0] n22995_o;
  wire n22997_o;
  wire [11:0] n22998_o;
  wire n23000_o;
  wire [11:0] n23001_o;
  wire n23003_o;
  wire [11:0] n23004_o;
  wire n23006_o;
  wire [11:0] n23007_o;
  wire [6:0] n23008_o;
  wire [11:0] n23009_o;
  reg [11:0] n23010_o;
  wire [11:0] n23011_o;
  reg [11:0] n23012_o;
  wire [11:0] n23013_o;
  reg [11:0] n23014_o;
  wire [11:0] n23015_o;
  reg [11:0] n23016_o;
  wire [11:0] n23017_o;
  reg [11:0] n23018_o;
  wire [11:0] n23019_o;
  reg [11:0] n23020_o;
  wire [11:0] n23021_o;
  reg [11:0] n23022_o;
  wire [11:0] n23023_o;
  reg [11:0] n23024_o;
  wire n23026_o;
  wire n23029_o;
  wire [95:0] n23030_o;
  wire [95:0] n23031_o;
  wire [95:0] n23032_o;
  wire [95:0] n23033_o;
  wire [95:0] n23034_o;
  wire n23036_o;
  wire [2:0] n23038_o;
  wire [2:0] n23040_o;
  wire n23045_o;
  wire [12:0] xregister_file_i_n23094;
  wire [255:0] xregister_file_i_n23095;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n23100;
  wire [12:0] iregister_i_n23101;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n23108_o;
  wire n23110_o;
  wire n23111_o;
  wire n23113_o;
  wire n23114_o;
  wire n23117_o;
  wire n23119_o;
  wire n23120_o;
  wire n23123_o;
  wire n23124_o;
  wire [4:0] n23132_o;
  wire n23133_o;
  wire [4:0] n23134_o;
  wire [4:0] n23137_o;
  wire [4:0] n23138_o;
  wire [4:0] n23139_o;
  wire n23140_o;
  wire n23141_o;
  wire n23142_o;
  wire n23143_o;
  wire n23144_o;
  wire n23145_o;
  wire n23146_o;
  wire n23147_o;
  wire n23148_o;
  wire n23151_o;
  wire [31:0] n23153_o;
  wire [11:0] n23154_o;
  wire [11:0] n23155_o;
  wire [31:0] alu_0_i_n23156;
  wire alu_0_i_n23157;
  wire [11:0] alu_0_i_n23158;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n23165_o;
  wire [11:0] n23166_o;
  wire [11:0] n23167_o;
  wire [31:0] alu_1_i_n23168;
  wire alu_1_i_n23169;
  wire [11:0] alu_1_i_n23170;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n23177_o;
  wire [11:0] n23178_o;
  wire [11:0] n23179_o;
  wire [31:0] alu_2_i_n23180;
  wire alu_2_i_n23181;
  wire [11:0] alu_2_i_n23182;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n23189_o;
  wire [11:0] n23190_o;
  wire [11:0] n23191_o;
  wire [31:0] alu_3_i_n23192;
  wire alu_3_i_n23193;
  wire [11:0] alu_3_i_n23194;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n23201_o;
  wire [11:0] n23202_o;
  wire [11:0] n23203_o;
  wire [31:0] alu_4_i_n23204;
  wire alu_4_i_n23205;
  wire [11:0] alu_4_i_n23206;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n23213_o;
  wire [11:0] n23214_o;
  wire [11:0] n23215_o;
  wire [31:0] alu_5_i_n23216;
  wire alu_5_i_n23217;
  wire [11:0] alu_5_i_n23218;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n23225_o;
  wire [11:0] n23226_o;
  wire [11:0] n23227_o;
  wire [31:0] alu_6_i_n23228;
  wire alu_6_i_n23229;
  wire [11:0] alu_6_i_n23230;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n23237_o;
  wire [11:0] n23238_o;
  wire [11:0] n23239_o;
  wire [31:0] alu_7_i_n23240;
  wire alu_7_i_n23241;
  wire [11:0] alu_7_i_n23242;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n23249_o;
  wire n23250_o;
  wire [12:0] ialu_i_n23251;
  wire ialu_i_n23252;
  wire ialu_i_n23253;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n23262;
  wire [95:0] register_bank_i_n23263;
  wire [16:0] n23264_o;
  wire [16:0] n23265_o;
  wire [95:0] register_bank_i_n23266;
  wire register_bank_i_n23267;
  wire register_bank_i_n23268;
  wire [2:0] register_bank_i_n23269;
  wire [2:0] register_bank_i_n23270;
  wire [1:0] register_bank_i_n23271;
  wire [2:0] register_bank_i_n23272;
  wire [2:0] register_bank_i_n23273;
  wire register_bank_i_n23274;
  wire [1:0] register_bank_i_n23275;
  wire [1:0] register_bank_i_n23276;
  wire register_bank_i_n23277;
  wire [1:0] register_bank_i_n23278;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n23311;
  wire instr_decoder2_i_n23312;
  wire [3:0] instr_decoder2_i_n23313;
  wire instr_decoder2_i_n23314;
  wire instr_decoder2_i_n23315;
  wire instr_decoder2_i_n23316;
  wire instr_decoder2_i_n23317;
  wire [11:0] instr_decoder2_i_n23318;
  wire [11:0] instr_decoder2_i_n23319;
  wire [11:0] instr_decoder2_i_n23320;
  wire instr_decoder2_i_n23321;
  wire instr_decoder2_i_n23322;
  wire instr_decoder2_i_n23323;
  wire [7:0] instr_decoder2_i_n23324;
  wire instr_decoder2_i_n23325;
  wire [11:0] instr_decoder2_i_n23326;
  wire instr_decoder2_i_n23327;
  wire instr_decoder2_i_n23328;
  wire [3:0] instr_decoder2_i_n23329;
  wire [3:0] instr_decoder2_i_n23330;
  wire instr_decoder2_i_n23331;
  wire instr_decoder2_i_n23332;
  wire [2:0] instr_decoder2_i_n23333;
  wire [12:0] instr_decoder2_i_n23334;
  wire instr_decoder2_i_n23335;
  wire [4:0] instr_decoder2_i_n23336;
  wire [12:0] instr_decoder2_i_n23337;
  wire [12:0] instr_decoder2_i_n23338;
  wire [7:0] instr_decoder2_i_n23339;
  wire [7:0] instr_decoder2_i_n23340;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n23401;
  wire instr_dispatch2_i1_n23402;
  wire [11:0] instr_dispatch2_i1_n23403;
  wire [11:0] instr_dispatch2_i1_n23404;
  wire instr_dispatch2_i1_n23405;
  wire instr_dispatch2_i1_n23406;
  wire instr_dispatch2_i1_n23407;
  wire instr_dispatch2_i1_n23408;
  wire instr_dispatch2_i1_n23409;
  wire instr_dispatch2_i1_n23410;
  wire instr_dispatch2_i1_n23411;
  wire instr_dispatch2_i1_n23412;
  wire [11:0] instr_dispatch2_i1_n23413;
  wire [7:0] instr_dispatch2_i1_n23414;
  wire [95:0] instr_dispatch2_i1_n23415;
  wire [7:0] instr_dispatch2_i1_n23416;
  wire [95:0] instr_dispatch2_i1_n23417;
  wire [95:0] instr_dispatch2_i1_n23418;
  wire [11:0] instr_dispatch2_i1_n23419;
  wire [4:0] instr_dispatch2_i1_n23420;
  wire [3:0] instr_dispatch2_i1_n23421;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n23467_o;
  wire [95:0] n23468_o;
  wire [7:0] n23469_o;
  wire [95:0] n23470_o;
  reg [95:0] n23471_q;
  wire [95:0] n23472_o;
  reg [95:0] n23473_q;
  reg n23474_q;
  reg n23475_q;
  wire n23476_o;
  reg n23477_q;
  wire [1:0] n23478_o;
  reg [1:0] n23479_q;
  wire [1:0] n23480_o;
  reg [1:0] n23481_q;
  wire [2:0] n23482_o;
  reg [2:0] n23483_q;
  wire [2:0] n23484_o;
  reg [2:0] n23485_q;
  wire n23486_o;
  reg n23487_q;
  wire [1:0] n23488_o;
  reg [1:0] n23489_q;
  reg [2:0] n23490_q;
  reg [2:0] n23491_q;
  reg [1:0] n23492_q;
  reg [2:0] n23495_q;
  reg [2:0] n23496_q;
  reg n23497_q;
  reg [1:0] n23498_q;
  reg [1:0] n23499_q;
  reg n23500_q;
  reg [1:0] n23501_q;
  reg [21:0] n23502_q;
  reg [2:0] n23503_q;
  reg [21:0] n23504_q;
  reg [95:0] n23505_q;
  wire n23506_o;
  reg n23507_q;
  wire n23508_o;
  reg n23509_q;
  wire n23510_o;
  reg n23511_q;
  wire n23512_o;
  reg n23513_q;
  reg [21:0] n23514_q;
  reg [21:0] n23515_q;
  wire [5:0] n23516_o;
  reg [5:0] n23517_q;
  wire n23518_o;
  reg n23519_q;
  wire [2:0] n23522_o;
  reg [2:0] n23523_q;
  wire [1:0] n23524_o;
  reg [1:0] n23525_q;
  wire n23526_o;
  reg n23527_q;
  wire [21:0] n23528_o;
  reg [21:0] n23529_q;
  wire n23530_o;
  reg n23531_q;
  wire [2:0] n23532_o;
  reg [2:0] n23533_q;
  wire [1:0] n23534_o;
  reg [1:0] n23535_q;
  wire n23536_o;
  wire n23537_o;
  wire n23538_o;
  reg n23539_q;
  wire n23540_o;
  wire n23541_o;
  wire [21:0] n23542_o;
  reg [21:0] n23543_q;
  wire n23544_o;
  reg n23545_q;
  wire [1:0] n23546_o;
  reg [1:0] n23547_q;
  wire [1:0] n23548_o;
  reg [1:0] n23549_q;
  wire n23550_o;
  reg n23551_q;
  wire [1:0] n23552_o;
  reg [1:0] n23553_q;
  reg [83:0] n23554_q;
  wire [95:0] n23555_o;
  reg [2:0] n23556_q;
  reg [2:0] n23557_q;
  reg [2:0] n23558_q;
  reg [79:0] n23560_q;
  reg [31:0] n23561_q;
  reg n23562_q;
  reg n23563_q;
  reg n23564_q;
  reg [1:0] n23565_q;
  reg [3:0] n23566_q;
  reg n23567_q;
  reg [3:0] n23568_q;
  reg n23569_q;
  reg [3:0] n23570_q;
  reg n23571_q;
  reg n23572_q;
  reg [1:0] n23573_q;
  reg [27:0] n23574_q;
  reg n23575_q;
  reg n23576_q;
  reg n23578_q;
  reg n23579_q;
  reg n23581_q;
  reg n23582_q;
  reg n23583_q;
  reg [21:0] n23584_q;
  reg n23585_q;
  reg [21:0] n23586_q;
  reg [21:0] n23587_q;
  reg n23588_q;
  reg [21:0] n23589_q;
  reg [5:0] n23590_q;
  reg n23591_q;
  reg n23592_q;
  reg n23593_q;
  reg [2:0] n23594_q;
  reg [1:0] n23595_q;
  reg n23596_q;
  reg n23597_q;
  reg [2:0] n23598_q;
  reg [1:0] n23599_q;
  reg n23600_q;
  reg [1:0] n23601_q;
  reg [1:0] n23602_q;
  reg n23603_q;
  reg [1:0] n23604_q;
  reg [95:0] n23605_q;
  reg n23606_q;
  wire [2:0] n23607_o;
  wire [2:0] n23608_o;
  assign i_y_neg_out = n23249_o;
  assign i_y_zero_out = n23250_o;
  assign dp_readdata_out = n22923_o;
  assign dp_readdata_vm_out = n22925_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n23607_o;
  assign dp_read_vaddr_out = n23608_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n22903_o;
  assign dp_read_data_type_out = n22905_o;
  assign dp_read_stream_out = n22907_o;
  assign dp_read_stream_id_out = n22909_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n23262; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n23263; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n23401; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n23402; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n23410; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n23407; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n23408; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n23409; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n23415; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n23416; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n23318; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n23319; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n23320; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n23101; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n23335; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n23311; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n23417; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n23418; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n23419; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n23467_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n23468_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n23469_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n23420; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n23421; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n23313; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n23151_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n23124_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n22917_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n23403; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n23404; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n23413; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n23414; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n22915_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n22916_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n23312; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n23317; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n23314; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n23315; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n23316; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n23325; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n23326; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n23321; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n23322; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n23323; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n23324; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n23405; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n23406; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n23412; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n23327; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n23328; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n23329; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n23100; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n23330; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n23331; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n23332; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n23333; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n23334; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n23471_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n23473_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n23474_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n23475_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n23477_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n23479_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n23481_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n23483_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n23485_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n23487_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n23489_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n23336; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n23337; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n23338; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n23251; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n23252; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n23253; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n23411; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n23339; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n23340; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n23094; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n23095; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n22583_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n22584_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n22623_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:191:8  */
  assign dp_wr_fork = n22624_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n22585_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n22625_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n22626_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n22627_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n22628_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n22629_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n22630_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n22631_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n22586_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n22587_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n22588_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n22589_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n22590_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n22591_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n22592_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n22593_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n22594_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n22595_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n22877_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n22596_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n22597_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n22633_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n22636_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n23490_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n23491_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n23492_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n23495_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n23496_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n23497_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n23498_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n23499_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n23500_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n23501_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n23502_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n23503_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n23504_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n23505_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n23507_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n23509_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n23511_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:238:8  */
  assign dp_wr_fork_r = n23513_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n23514_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n23515_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n23517_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n23519_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n23523_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n23525_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n23527_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n23529_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n23531_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n23533_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n23535_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n23539_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n23543_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n23545_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n23547_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n23549_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n23551_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n23553_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n23555_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n23556_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n23557_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n23558_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n22901_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n22562_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n23268; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n23269; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n23270; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n23271; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n23272; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n23273; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n23266; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n23267; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n23274; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n23275; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n23276; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n23277; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n23278; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n22440_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n22441_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n22442_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n23560_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n23561_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n23562_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n23563_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n23564_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n23565_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n23566_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n23567_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n23568_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n23569_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n23570_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n23571_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n23572_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n23573_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n23574_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n23575_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n23576_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n23578_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n23579_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n23581_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n23582_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n23583_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n23584_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n23585_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n23586_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n23587_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n23588_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n23589_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n23590_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n23591_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n23592_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n23593_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n23594_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n23595_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n23596_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n23597_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n23598_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n23599_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n23600_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n23601_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n23602_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n23603_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n23604_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n23605_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n23606_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n22440_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n22441_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n22442_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n22445_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n22533_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n22534_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n22535_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n22536_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n22539_o = n22536_o ? 3'b001 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n22541_o = n22535_o + n22533_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n22542_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n22543_o = n22542_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n22544_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n22545_o = n22544_o & n22543_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n22546_o = n22533_o & n22535_o;
  /* ../../HW/src/pcore/pcore.vhd:104:8  */
  assign n22547_o = {n22539_o, 2'b01};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n22548_o = n22533_o & n22547_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n22549_o = n22546_o == n22548_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n22550_o = n22549_o & n22534_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n22551_o = ~n22534_o;
  /* ../../HW/src/pcore/pcore.vhd:349:1  */
  assign n22552_o = {n22539_o, 2'b01};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n22553_o = $unsigned(n22552_o) >= $unsigned(n22535_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n22554_o = n22553_o & n22551_o;
  /* ../../HW/src/pcore/pcore.vhd:349:1  */
  assign n22555_o = {n22539_o, 2'b01};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n22556_o = $unsigned(n22555_o) <= $unsigned(n22541_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n22557_o = n22556_o & n22554_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n22558_o = n22550_o | n22557_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n22559_o = n22558_o & n22545_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n22562_o = n22559_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n22568_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n22570_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n22572_o = n22570_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n22574_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n22575_o = n22574_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n22576_o = dp_read_gen_valid_in_r & n22575_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n22578_o = n22576_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n22580_o = n22576_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n22582_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22583_o = n22568_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22584_o = n22568_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22585_o = n22568_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22586_o = n22568_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22587_o = n22568_o ? n22572_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22588_o = n22568_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22589_o = n22568_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22590_o = n22568_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22591_o = n22568_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22592_o = n22568_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22593_o = n22568_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22594_o = n22568_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22595_o = n22568_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22596_o = n22568_o ? n22578_o : n22582_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n22597_o = n22568_o ? n22580_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n22602_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n22603_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n22604_o = dp_write_in_r & n22603_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n22605_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n22606_o = n22604_o & n22605_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n22608_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n22610_o = n22608_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n22612_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n22613_o = n22612_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n22614_o = dp_write_gen_valid_in_r & n22613_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n22616_o = n22614_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n22620_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n22622_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22623_o = n22602_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22624_o = n22602_o ? dp_wr_fork_in_r : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22625_o = n22602_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22626_o = n22602_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22627_o = n22602_o ? n22606_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22628_o = n22602_o ? n22610_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22629_o = n22602_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22630_o = n22602_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22631_o = n22602_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22633_o = n22602_o ? n22616_o : n22620_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n22636_o = n22602_o ? 3'b000 : n22622_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n22641_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n22644_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n22645_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n22646_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n22648_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n22649_o = n22645_o ? n22646_o : n22648_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n22651_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n22652_o = n22644_o ? n22649_o : n22651_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n22654_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n22718_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n22787_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n22790_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n22791_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n22792_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n22794_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n22795_o = n22791_o ? n22792_o : n22794_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n22797_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n22798_o = n22790_o ? n22795_o : n22797_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n22800_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n22801_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n22802_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n22812_o = n22800_o ? n22801_o : n22802_o;
  assign n22854_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n22855_o = n22787_o ? 12'b000000000000 : n22854_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n22869_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n22871_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n22872_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n22873_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n22874_o = n22871_o ? n22872_o : n22873_o;
  assign n22876_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n22874_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n22877_o = n22869_o ? n22876_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n22883_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n22884_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n22885_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n22887_o = n22883_o == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n22888_o = n22887_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n22890_o = n22884_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n22891_o = n22890_o & n22888_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n22894_o = n22891_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n22896_o = n22883_o == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n22897_o = n22896_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n22900_o = n22897_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n22901_o = n22885_o ? n22894_o : n22900_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n22903_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n22905_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n22907_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n22909_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n22915_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n22916_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n22917_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n22920_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n22921_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n22923_o = n22920_o ? 96'bZ : n22921_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n22925_o = n22920_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n22930_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n22981_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n22984_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n22985_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n22986_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n22988_o = n22985_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n22989_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n22991_o = n22985_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n22992_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n22994_o = n22985_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n22995_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n22997_o = n22985_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n22998_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n23000_o = n22985_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n23001_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n23003_o = n22985_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n23004_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n23006_o = n22985_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n23007_o = dp_readdata_vm[11:0];
  assign n23008_o = {n23006_o, n23003_o, n23000_o, n22997_o, n22994_o, n22991_o, n22988_o};
  assign n23009_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23010_o = n23009_o;
      7'b0100000: n23010_o = n23009_o;
      7'b0010000: n23010_o = n23009_o;
      7'b0001000: n23010_o = n23009_o;
      7'b0000100: n23010_o = n23009_o;
      7'b0000010: n23010_o = n23009_o;
      7'b0000001: n23010_o = n23009_o;
      default: n23010_o = n23007_o;
    endcase
  assign n23011_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23012_o = n23004_o;
      7'b0100000: n23012_o = n23011_o;
      7'b0010000: n23012_o = n23011_o;
      7'b0001000: n23012_o = n23011_o;
      7'b0000100: n23012_o = n23011_o;
      7'b0000010: n23012_o = n23011_o;
      7'b0000001: n23012_o = n23011_o;
      default: n23012_o = n23011_o;
    endcase
  assign n23013_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23014_o = n23013_o;
      7'b0100000: n23014_o = n23001_o;
      7'b0010000: n23014_o = n23013_o;
      7'b0001000: n23014_o = n23013_o;
      7'b0000100: n23014_o = n23013_o;
      7'b0000010: n23014_o = n23013_o;
      7'b0000001: n23014_o = n23013_o;
      default: n23014_o = n23013_o;
    endcase
  assign n23015_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23016_o = n23015_o;
      7'b0100000: n23016_o = n23015_o;
      7'b0010000: n23016_o = n22998_o;
      7'b0001000: n23016_o = n23015_o;
      7'b0000100: n23016_o = n23015_o;
      7'b0000010: n23016_o = n23015_o;
      7'b0000001: n23016_o = n23015_o;
      default: n23016_o = n23015_o;
    endcase
  assign n23017_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23018_o = n23017_o;
      7'b0100000: n23018_o = n23017_o;
      7'b0010000: n23018_o = n23017_o;
      7'b0001000: n23018_o = n22995_o;
      7'b0000100: n23018_o = n23017_o;
      7'b0000010: n23018_o = n23017_o;
      7'b0000001: n23018_o = n23017_o;
      default: n23018_o = n23017_o;
    endcase
  assign n23019_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23020_o = n23019_o;
      7'b0100000: n23020_o = n23019_o;
      7'b0010000: n23020_o = n23019_o;
      7'b0001000: n23020_o = n23019_o;
      7'b0000100: n23020_o = n22992_o;
      7'b0000010: n23020_o = n23019_o;
      7'b0000001: n23020_o = n23019_o;
      default: n23020_o = n23019_o;
    endcase
  assign n23021_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23022_o = n23021_o;
      7'b0100000: n23022_o = n23021_o;
      7'b0010000: n23022_o = n23021_o;
      7'b0001000: n23022_o = n23021_o;
      7'b0000100: n23022_o = n23021_o;
      7'b0000010: n23022_o = n22989_o;
      7'b0000001: n23022_o = n23021_o;
      default: n23022_o = n23021_o;
    endcase
  assign n23023_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n23008_o)
      7'b1000000: n23024_o = n23023_o;
      7'b0100000: n23024_o = n23023_o;
      7'b0010000: n23024_o = n23023_o;
      7'b0001000: n23024_o = n23023_o;
      7'b0000100: n23024_o = n23023_o;
      7'b0000010: n23024_o = n23023_o;
      7'b0000001: n23024_o = n22986_o;
      default: n23024_o = n23023_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n23026_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n23029_o = n23026_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n23030_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n23031_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n23032_o = {n23024_o, n23022_o, n23020_o, n23018_o, n23016_o, n23014_o, n23012_o, n23010_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n23033_o = n22984_o ? n23032_o : n23030_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n23034_o = n22984_o ? dp_readdata2_r : n23031_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n23036_o = n22984_o ? n23029_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n23038_o = n22984_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n23040_o = n22984_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n23045_o = dp_readena_vm ? n23036_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n23094 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n23095 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n23100 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n23101 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n23108_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n23110_o = dp_rd_pid == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n23111_o = n23110_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n23113_o = dp_rd_cid == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n23114_o = n23113_o & n23111_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n23117_o = n23114_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n23119_o = dp_rd_pid == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n23120_o = n23119_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n23123_o = n23120_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n23124_o = n23108_o ? n23117_o : n23123_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n23132_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n23133_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n23134_o = dp_mcast_addr + n23132_o;
  /* ../../HW/src/pcore/pcore.vhd:1022:1  */
  assign n23137_o = dp_wr_fork ? 5'b00001 : 5'b00101;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n23138_o = n23132_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n23139_o = n23132_o & n23137_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n23140_o = n23138_o == n23139_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n23141_o = n23140_o & n23133_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n23142_o = ~n23133_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n23143_o = $unsigned(n23137_o) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n23144_o = n23143_o & n23142_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n23145_o = $unsigned(n23137_o) <= $unsigned(n23134_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n23146_o = n23145_o & n23144_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n23147_o = n23141_o | n23146_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n23148_o = n23147_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n23151_o = n23148_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n23153_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n23154_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n23155_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n23156 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n23157 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n23158 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23153_o),
    .x1_in(n23154_o),
    .x2_in(n23155_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n23165_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n23166_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n23167_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n23168 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n23169 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n23170 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23165_o),
    .x1_in(n23166_o),
    .x2_in(n23167_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n23177_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n23178_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n23179_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n23180 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n23181 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n23182 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23177_o),
    .x1_in(n23178_o),
    .x2_in(n23179_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n23189_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n23190_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n23191_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n23192 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n23193 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n23194 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23189_o),
    .x1_in(n23190_o),
    .x2_in(n23191_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n23201_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n23202_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n23203_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n23204 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n23205 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n23206 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23201_o),
    .x1_in(n23202_o),
    .x2_in(n23203_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n23213_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n23214_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n23215_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n23216 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n23217 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n23218 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23213_o),
    .x1_in(n23214_o),
    .x2_in(n23215_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n23225_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n23226_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n23227_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n23228 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n23229 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n23230 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23225_o),
    .x1_in(n23226_o),
    .x2_in(n23227_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n23237_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n23238_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n23239_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n23240 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n23241 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n23242 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n23237_o),
    .x1_in(n23238_o),
    .x2_in(n23239_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n23249_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n23250_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n23251 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n23252 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n23253 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n23262 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n23263 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n23264_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n23265_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n23266 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n23267 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n23268 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n23269 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n23270 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n23271 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n23272 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n23273 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n23274 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n23275 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n23276 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n23277 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n23278 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n23264_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n23265_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n23311 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n23312 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n23313 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n23314 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n23315 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n23316 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n23317 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n23318 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n23319 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n23320 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n23321 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n23322 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n23323 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n23324 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n23325 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n23326 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n23327 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n23328 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n23329 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n23330 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n23331 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n23332 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n23333 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n23334 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n23335 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n23336 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n23337 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n23338 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n23339 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n23340 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_1_1 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n23401 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n23402 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n23403 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n23404 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n23405 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n23406 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n23407 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n23408 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n23409 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n23410 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n23411 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n23412 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n23413 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n23414 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n23415 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n23416 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n23417 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n23418 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n23419 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n23420 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n23421 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n23467_o = {alu_7_i_n23240, alu_6_i_n23228, alu_5_i_n23216, alu_4_i_n23204, alu_3_i_n23192, alu_2_i_n23180, alu_1_i_n23168, alu_0_i_n23156};
  assign n23468_o = {alu_7_i_n23242, alu_6_i_n23230, alu_5_i_n23218, alu_4_i_n23206, alu_3_i_n23194, alu_2_i_n23182, alu_1_i_n23170, alu_0_i_n23158};
  assign n23469_o = {alu_7_i_n23241, alu_6_i_n23229, alu_5_i_n23217, alu_4_i_n23205, alu_3_i_n23193, alu_2_i_n23181, alu_1_i_n23169, alu_0_i_n23157};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23470_o = dp_readena_vm ? n23033_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23471_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n23471_q <= n23470_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23472_o = dp_readena_vm ? n23034_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23473_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n23473_q <= n23472_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23474_q <= 1'b0;
    else
      n23474_q <= n23045_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23475_q <= 1'b0;
    else
      n23475_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23476_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23477_q <= 1'b0;
    else
      n23477_q <= n23476_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23478_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23479_q <= 2'b00;
    else
      n23479_q <= n23478_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23480_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23481_q <= 2'b00;
    else
      n23481_q <= n23480_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23482_o = dp_readena_vm ? n23038_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23483_q <= 3'b000;
    else
      n23483_q <= n23482_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23484_o = dp_readena_vm ? n23040_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23485_q <= 3'b000;
    else
      n23485_q <= n23484_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23486_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23487_q <= 1'b0;
    else
      n23487_q <= n23486_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n23488_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n22981_o)
    if (n22981_o)
      n23489_q <= 2'b00;
    else
      n23489_q <= n23488_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23490_q <= 3'b000;
    else
      n23490_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23491_q <= 3'b000;
    else
      n23491_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23492_q <= 2'b00;
    else
      n23492_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23495_q <= 3'b000;
    else
      n23495_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23496_q <= 3'b000;
    else
      n23496_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23497_q <= 1'b0;
    else
      n23497_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23498_q <= 2'b00;
    else
      n23498_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23499_q <= 2'b00;
    else
      n23499_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23500_q <= 1'b0;
    else
      n23500_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23501_q <= 2'b00;
    else
      n23501_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23502_q <= 22'b0000000000000000000000;
    else
      n23502_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23503_q <= 3'b000;
    else
      n23503_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23504_q <= 22'b0000000000000000000000;
    else
      n23504_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23505_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n23505_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23506_o = n22654_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23507_q <= 1'b0;
    else
      n23507_q <= n23506_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23508_o = n22654_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23509_q <= 1'b0;
    else
      n23509_q <= n23508_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23510_o = n22800_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23511_q <= 1'b0;
    else
      n23511_q <= n23510_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23512_o = n22800_o ? dp_wr_fork : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23513_q <= 1'b0;
    else
      n23513_q <= n23512_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23514_q <= 22'b0000000000000000000000;
    else
      n23514_q <= n22652_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23515_q <= 22'b0000000000000000000000;
    else
      n23515_q <= n22798_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23516_o = n22800_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23517_q <= 6'b000000;
    else
      n23517_q <= n23516_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23518_o = n22800_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23519_q <= 1'b0;
    else
      n23519_q <= n23518_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23522_o = n22800_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23523_q <= 3'b000;
    else
      n23523_q <= n23522_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23524_o = n22800_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23525_q <= 2'b00;
    else
      n23525_q <= n23524_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23526_o = n22800_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23527_q <= 1'b0;
    else
      n23527_q <= n23526_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n23528_o = n22800_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23529_q <= 22'b0000000000000000000000;
    else
      n23529_q <= n23528_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23530_o = n22654_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23531_q <= 1'b0;
    else
      n23531_q <= n23530_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23532_o = n22654_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23533_q <= 3'b000;
    else
      n23533_q <= n23532_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23534_o = n22654_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23535_q <= 2'b00;
    else
      n23535_q <= n23534_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n23536_o = ~n22641_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n23537_o = n22654_o & n23536_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23538_o = n23537_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n23539_q <= n23538_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n23540_o = ~n22641_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n23541_o = n22654_o & n23540_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23542_o = n23541_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n23543_q <= n23542_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23544_o = n22654_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23545_q <= 1'b0;
    else
      n23545_q <= n23544_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23546_o = n22654_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23547_q <= 2'b00;
    else
      n23547_q <= n23546_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23548_o = n22654_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23549_q <= 2'b00;
    else
      n23549_q <= n23548_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23550_o = n22654_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23551_q <= 1'b0;
    else
      n23551_q <= n23550_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n23552_o = n22654_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23553_q <= 2'b00;
    else
      n23553_q <= n23552_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23554_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n23554_q <= n22812_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n23555_o = {n22855_o, n23554_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23556_q <= 3'b000;
    else
      n23556_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n22641_o)
    if (n22641_o)
      n23557_q <= 3'b000;
    else
      n23557_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n22787_o)
    if (n22787_o)
      n23558_q <= 3'b000;
    else
      n23558_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23560_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n23560_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23561_q <= 32'b00000000000000000000000000000000;
    else
      n23561_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23562_q <= 1'b0;
    else
      n23562_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23563_q <= 1'b0;
    else
      n23563_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23564_q <= 1'b0;
    else
      n23564_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23565_q <= 2'b00;
    else
      n23565_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23566_q <= 4'b0000;
    else
      n23566_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23567_q <= 1'b0;
    else
      n23567_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23568_q <= 4'b0000;
    else
      n23568_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23569_q <= 1'b0;
    else
      n23569_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23570_q <= 4'b0000;
    else
      n23570_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23571_q <= 1'b0;
    else
      n23571_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23572_q <= 1'b0;
    else
      n23572_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23573_q <= 2'b00;
    else
      n23573_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n22930_o)
    if (n22930_o)
      n23574_q <= 28'b0000000000000000000000000000;
    else
      n23574_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23575_q <= 1'b0;
    else
      n23575_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23576_q <= 1'b0;
    else
      n23576_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23578_q <= 1'b0;
    else
      n23578_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n22718_o)
    if (n22718_o)
      n23579_q <= 1'b0;
    else
      n23579_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23581_q <= 1'b0;
    else
      n23581_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23582_q <= 1'b0;
    else
      n23582_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23583_q <= 1'b0;
    else
      n23583_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23584_q <= 22'b0000000000000000000000;
    else
      n23584_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23585_q <= 1'b0;
    else
      n23585_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23586_q <= 22'b0000000000000000000000;
    else
      n23586_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23587_q <= 22'b0000000000000000000000;
    else
      n23587_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23588_q <= 1'b0;
    else
      n23588_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23589_q <= 22'b0000000000000000000000;
    else
      n23589_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23590_q <= 6'b000000;
    else
      n23590_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23591_q <= 1'b0;
    else
      n23591_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23592_q <= 1'b0;
    else
      n23592_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23593_q <= 1'b0;
    else
      n23593_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23594_q <= 3'b000;
    else
      n23594_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23595_q <= 2'b00;
    else
      n23595_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23596_q <= 1'b0;
    else
      n23596_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23597_q <= 1'b0;
    else
      n23597_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23598_q <= 3'b000;
    else
      n23598_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23599_q <= 2'b00;
    else
      n23599_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23600_q <= 1'b0;
    else
      n23600_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23601_q <= 2'b00;
    else
      n23601_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23602_q <= 2'b00;
    else
      n23602_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23603_q <= 1'b0;
    else
      n23603_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23604_q <= 2'b00;
    else
      n23604_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23605_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n23605_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n22445_o)
    if (n22445_o)
      n23606_q <= 1'b0;
    else
      n23606_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n23607_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n23608_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_1_0
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire dp_wr_fork;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire dp_wr_fork_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n21259_o;
  wire n21260_o;
  wire n21261_o;
  wire n21264_o;
  wire [4:0] n21352_o;
  wire n21353_o;
  wire [4:0] n21354_o;
  wire n21355_o;
  wire [2:0] n21358_o;
  wire [4:0] n21360_o;
  wire n21361_o;
  wire n21362_o;
  wire n21363_o;
  wire n21364_o;
  wire [4:0] n21365_o;
  wire [4:0] n21366_o;
  wire [4:0] n21367_o;
  wire n21368_o;
  wire n21369_o;
  wire n21370_o;
  wire [4:0] n21371_o;
  wire n21372_o;
  wire n21373_o;
  wire [4:0] n21374_o;
  wire n21375_o;
  wire n21376_o;
  wire n21377_o;
  wire n21378_o;
  wire n21381_o;
  wire n21387_o;
  wire n21389_o;
  wire [2:0] n21391_o;
  wire n21393_o;
  wire n21394_o;
  wire n21395_o;
  wire [2:0] n21397_o;
  wire [2:0] n21399_o;
  wire [2:0] n21401_o;
  wire n21402_o;
  wire n21403_o;
  wire [21:0] n21404_o;
  wire n21405_o;
  wire [2:0] n21406_o;
  wire [1:0] n21407_o;
  wire n21408_o;
  wire [21:0] n21409_o;
  wire n21410_o;
  wire [1:0] n21411_o;
  wire [1:0] n21412_o;
  wire n21413_o;
  wire [1:0] n21414_o;
  wire [2:0] n21415_o;
  wire [2:0] n21416_o;
  wire n21421_o;
  wire n21422_o;
  wire n21423_o;
  wire n21424_o;
  wire n21425_o;
  wire n21427_o;
  wire [2:0] n21429_o;
  wire n21431_o;
  wire n21432_o;
  wire n21433_o;
  wire [2:0] n21435_o;
  wire [2:0] n21439_o;
  wire [2:0] n21441_o;
  wire n21442_o;
  wire n21443_o;
  wire [21:0] n21444_o;
  wire [5:0] n21445_o;
  wire n21446_o;
  wire [2:0] n21447_o;
  wire [1:0] n21448_o;
  wire n21449_o;
  wire [21:0] n21450_o;
  wire [2:0] n21452_o;
  wire [2:0] n21455_o;
  wire n21460_o;
  wire n21463_o;
  wire n21464_o;
  wire [21:0] n21465_o;
  wire [21:0] n21467_o;
  wire [21:0] n21468_o;
  wire [21:0] n21470_o;
  wire [21:0] n21471_o;
  wire n21473_o;
  wire n21537_o;
  wire n21606_o;
  wire n21609_o;
  wire n21610_o;
  wire [21:0] n21611_o;
  wire [21:0] n21613_o;
  wire [21:0] n21614_o;
  wire [21:0] n21616_o;
  wire [21:0] n21617_o;
  wire n21619_o;
  wire [83:0] n21620_o;
  wire [83:0] n21621_o;
  wire [83:0] n21631_o;
  wire [11:0] n21673_o;
  wire [11:0] n21674_o;
  wire n21688_o;
  wire n21690_o;
  wire [11:0] n21691_o;
  wire [11:0] n21692_o;
  wire [11:0] n21693_o;
  wire [95:0] n21695_o;
  wire [95:0] n21696_o;
  wire [1:0] n21702_o;
  wire [2:0] n21703_o;
  wire n21704_o;
  wire n21706_o;
  wire n21707_o;
  wire n21709_o;
  wire n21710_o;
  wire n21713_o;
  wire n21715_o;
  wire n21716_o;
  wire n21719_o;
  wire n21720_o;
  wire [1:0] n21722_o;
  wire [1:0] n21724_o;
  wire n21726_o;
  wire [1:0] n21728_o;
  wire [1:0] n21734_o;
  wire [2:0] n21735_o;
  wire [4:0] n21736_o;
  wire n21739_o;
  wire [95:0] n21740_o;
  wire [95:0] n21742_o;
  wire n21744_o;
  wire n21749_o;
  wire n21800_o;
  wire n21803_o;
  wire [2:0] n21804_o;
  wire [11:0] n21805_o;
  wire n21807_o;
  wire [11:0] n21808_o;
  wire n21810_o;
  wire [11:0] n21811_o;
  wire n21813_o;
  wire [11:0] n21814_o;
  wire n21816_o;
  wire [11:0] n21817_o;
  wire n21819_o;
  wire [11:0] n21820_o;
  wire n21822_o;
  wire [11:0] n21823_o;
  wire n21825_o;
  wire [11:0] n21826_o;
  wire [6:0] n21827_o;
  wire [11:0] n21828_o;
  reg [11:0] n21829_o;
  wire [11:0] n21830_o;
  reg [11:0] n21831_o;
  wire [11:0] n21832_o;
  reg [11:0] n21833_o;
  wire [11:0] n21834_o;
  reg [11:0] n21835_o;
  wire [11:0] n21836_o;
  reg [11:0] n21837_o;
  wire [11:0] n21838_o;
  reg [11:0] n21839_o;
  wire [11:0] n21840_o;
  reg [11:0] n21841_o;
  wire [11:0] n21842_o;
  reg [11:0] n21843_o;
  wire n21845_o;
  wire n21848_o;
  wire [95:0] n21849_o;
  wire [95:0] n21850_o;
  wire [95:0] n21851_o;
  wire [95:0] n21852_o;
  wire [95:0] n21853_o;
  wire n21855_o;
  wire [2:0] n21857_o;
  wire [2:0] n21859_o;
  wire n21864_o;
  wire [12:0] xregister_file_i_n21913;
  wire [255:0] xregister_file_i_n21914;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n21919;
  wire [12:0] iregister_i_n21920;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n21927_o;
  wire n21929_o;
  wire n21930_o;
  wire n21932_o;
  wire n21933_o;
  wire n21936_o;
  wire n21938_o;
  wire n21939_o;
  wire n21942_o;
  wire n21943_o;
  wire [4:0] n21951_o;
  wire n21952_o;
  wire [4:0] n21953_o;
  wire [4:0] n21956_o;
  wire [4:0] n21957_o;
  wire [4:0] n21958_o;
  wire n21959_o;
  wire n21960_o;
  wire n21961_o;
  wire n21962_o;
  wire n21963_o;
  wire n21964_o;
  wire n21965_o;
  wire n21966_o;
  wire n21967_o;
  wire n21970_o;
  wire [31:0] n21972_o;
  wire [11:0] n21973_o;
  wire [11:0] n21974_o;
  wire [31:0] alu_0_i_n21975;
  wire alu_0_i_n21976;
  wire [11:0] alu_0_i_n21977;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n21984_o;
  wire [11:0] n21985_o;
  wire [11:0] n21986_o;
  wire [31:0] alu_1_i_n21987;
  wire alu_1_i_n21988;
  wire [11:0] alu_1_i_n21989;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n21996_o;
  wire [11:0] n21997_o;
  wire [11:0] n21998_o;
  wire [31:0] alu_2_i_n21999;
  wire alu_2_i_n22000;
  wire [11:0] alu_2_i_n22001;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n22008_o;
  wire [11:0] n22009_o;
  wire [11:0] n22010_o;
  wire [31:0] alu_3_i_n22011;
  wire alu_3_i_n22012;
  wire [11:0] alu_3_i_n22013;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n22020_o;
  wire [11:0] n22021_o;
  wire [11:0] n22022_o;
  wire [31:0] alu_4_i_n22023;
  wire alu_4_i_n22024;
  wire [11:0] alu_4_i_n22025;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n22032_o;
  wire [11:0] n22033_o;
  wire [11:0] n22034_o;
  wire [31:0] alu_5_i_n22035;
  wire alu_5_i_n22036;
  wire [11:0] alu_5_i_n22037;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n22044_o;
  wire [11:0] n22045_o;
  wire [11:0] n22046_o;
  wire [31:0] alu_6_i_n22047;
  wire alu_6_i_n22048;
  wire [11:0] alu_6_i_n22049;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n22056_o;
  wire [11:0] n22057_o;
  wire [11:0] n22058_o;
  wire [31:0] alu_7_i_n22059;
  wire alu_7_i_n22060;
  wire [11:0] alu_7_i_n22061;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n22068_o;
  wire n22069_o;
  wire [12:0] ialu_i_n22070;
  wire ialu_i_n22071;
  wire ialu_i_n22072;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n22081;
  wire [95:0] register_bank_i_n22082;
  wire [16:0] n22083_o;
  wire [16:0] n22084_o;
  wire [95:0] register_bank_i_n22085;
  wire register_bank_i_n22086;
  wire register_bank_i_n22087;
  wire [2:0] register_bank_i_n22088;
  wire [2:0] register_bank_i_n22089;
  wire [1:0] register_bank_i_n22090;
  wire [2:0] register_bank_i_n22091;
  wire [2:0] register_bank_i_n22092;
  wire register_bank_i_n22093;
  wire [1:0] register_bank_i_n22094;
  wire [1:0] register_bank_i_n22095;
  wire register_bank_i_n22096;
  wire [1:0] register_bank_i_n22097;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n22130;
  wire instr_decoder2_i_n22131;
  wire [3:0] instr_decoder2_i_n22132;
  wire instr_decoder2_i_n22133;
  wire instr_decoder2_i_n22134;
  wire instr_decoder2_i_n22135;
  wire instr_decoder2_i_n22136;
  wire [11:0] instr_decoder2_i_n22137;
  wire [11:0] instr_decoder2_i_n22138;
  wire [11:0] instr_decoder2_i_n22139;
  wire instr_decoder2_i_n22140;
  wire instr_decoder2_i_n22141;
  wire instr_decoder2_i_n22142;
  wire [7:0] instr_decoder2_i_n22143;
  wire instr_decoder2_i_n22144;
  wire [11:0] instr_decoder2_i_n22145;
  wire instr_decoder2_i_n22146;
  wire instr_decoder2_i_n22147;
  wire [3:0] instr_decoder2_i_n22148;
  wire [3:0] instr_decoder2_i_n22149;
  wire instr_decoder2_i_n22150;
  wire instr_decoder2_i_n22151;
  wire [2:0] instr_decoder2_i_n22152;
  wire [12:0] instr_decoder2_i_n22153;
  wire instr_decoder2_i_n22154;
  wire [4:0] instr_decoder2_i_n22155;
  wire [12:0] instr_decoder2_i_n22156;
  wire [12:0] instr_decoder2_i_n22157;
  wire [7:0] instr_decoder2_i_n22158;
  wire [7:0] instr_decoder2_i_n22159;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n22220;
  wire instr_dispatch2_i1_n22221;
  wire [11:0] instr_dispatch2_i1_n22222;
  wire [11:0] instr_dispatch2_i1_n22223;
  wire instr_dispatch2_i1_n22224;
  wire instr_dispatch2_i1_n22225;
  wire instr_dispatch2_i1_n22226;
  wire instr_dispatch2_i1_n22227;
  wire instr_dispatch2_i1_n22228;
  wire instr_dispatch2_i1_n22229;
  wire instr_dispatch2_i1_n22230;
  wire instr_dispatch2_i1_n22231;
  wire [11:0] instr_dispatch2_i1_n22232;
  wire [7:0] instr_dispatch2_i1_n22233;
  wire [95:0] instr_dispatch2_i1_n22234;
  wire [7:0] instr_dispatch2_i1_n22235;
  wire [95:0] instr_dispatch2_i1_n22236;
  wire [95:0] instr_dispatch2_i1_n22237;
  wire [11:0] instr_dispatch2_i1_n22238;
  wire [4:0] instr_dispatch2_i1_n22239;
  wire [3:0] instr_dispatch2_i1_n22240;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n22286_o;
  wire [95:0] n22287_o;
  wire [7:0] n22288_o;
  wire [95:0] n22289_o;
  reg [95:0] n22290_q;
  wire [95:0] n22291_o;
  reg [95:0] n22292_q;
  reg n22293_q;
  reg n22294_q;
  wire n22295_o;
  reg n22296_q;
  wire [1:0] n22297_o;
  reg [1:0] n22298_q;
  wire [1:0] n22299_o;
  reg [1:0] n22300_q;
  wire [2:0] n22301_o;
  reg [2:0] n22302_q;
  wire [2:0] n22303_o;
  reg [2:0] n22304_q;
  wire n22305_o;
  reg n22306_q;
  wire [1:0] n22307_o;
  reg [1:0] n22308_q;
  reg [2:0] n22309_q;
  reg [2:0] n22310_q;
  reg [1:0] n22311_q;
  reg [2:0] n22314_q;
  reg [2:0] n22315_q;
  reg n22316_q;
  reg [1:0] n22317_q;
  reg [1:0] n22318_q;
  reg n22319_q;
  reg [1:0] n22320_q;
  reg [21:0] n22321_q;
  reg [2:0] n22322_q;
  reg [21:0] n22323_q;
  reg [95:0] n22324_q;
  wire n22325_o;
  reg n22326_q;
  wire n22327_o;
  reg n22328_q;
  wire n22329_o;
  reg n22330_q;
  wire n22331_o;
  reg n22332_q;
  reg [21:0] n22333_q;
  reg [21:0] n22334_q;
  wire [5:0] n22335_o;
  reg [5:0] n22336_q;
  wire n22337_o;
  reg n22338_q;
  wire [2:0] n22341_o;
  reg [2:0] n22342_q;
  wire [1:0] n22343_o;
  reg [1:0] n22344_q;
  wire n22345_o;
  reg n22346_q;
  wire [21:0] n22347_o;
  reg [21:0] n22348_q;
  wire n22349_o;
  reg n22350_q;
  wire [2:0] n22351_o;
  reg [2:0] n22352_q;
  wire [1:0] n22353_o;
  reg [1:0] n22354_q;
  wire n22355_o;
  wire n22356_o;
  wire n22357_o;
  reg n22358_q;
  wire n22359_o;
  wire n22360_o;
  wire [21:0] n22361_o;
  reg [21:0] n22362_q;
  wire n22363_o;
  reg n22364_q;
  wire [1:0] n22365_o;
  reg [1:0] n22366_q;
  wire [1:0] n22367_o;
  reg [1:0] n22368_q;
  wire n22369_o;
  reg n22370_q;
  wire [1:0] n22371_o;
  reg [1:0] n22372_q;
  reg [83:0] n22373_q;
  wire [95:0] n22374_o;
  reg [2:0] n22375_q;
  reg [2:0] n22376_q;
  reg [2:0] n22377_q;
  reg [79:0] n22379_q;
  reg [31:0] n22380_q;
  reg n22381_q;
  reg n22382_q;
  reg n22383_q;
  reg [1:0] n22384_q;
  reg [3:0] n22385_q;
  reg n22386_q;
  reg [3:0] n22387_q;
  reg n22388_q;
  reg [3:0] n22389_q;
  reg n22390_q;
  reg n22391_q;
  reg [1:0] n22392_q;
  reg [27:0] n22393_q;
  reg n22394_q;
  reg n22395_q;
  reg n22397_q;
  reg n22398_q;
  reg n22400_q;
  reg n22401_q;
  reg n22402_q;
  reg [21:0] n22403_q;
  reg n22404_q;
  reg [21:0] n22405_q;
  reg [21:0] n22406_q;
  reg n22407_q;
  reg [21:0] n22408_q;
  reg [5:0] n22409_q;
  reg n22410_q;
  reg n22411_q;
  reg n22412_q;
  reg [2:0] n22413_q;
  reg [1:0] n22414_q;
  reg n22415_q;
  reg n22416_q;
  reg [2:0] n22417_q;
  reg [1:0] n22418_q;
  reg n22419_q;
  reg [1:0] n22420_q;
  reg [1:0] n22421_q;
  reg n22422_q;
  reg [1:0] n22423_q;
  reg [95:0] n22424_q;
  reg n22425_q;
  wire [2:0] n22426_o;
  wire [2:0] n22427_o;
  assign i_y_neg_out = n22068_o;
  assign i_y_zero_out = n22069_o;
  assign dp_readdata_out = n21742_o;
  assign dp_readdata_vm_out = n21744_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n22426_o;
  assign dp_read_vaddr_out = n22427_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n21722_o;
  assign dp_read_data_type_out = n21724_o;
  assign dp_read_stream_out = n21726_o;
  assign dp_read_stream_id_out = n21728_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n22081; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n22082; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n22220; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n22221; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n22229; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n22226; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n22227; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n22228; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n22234; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n22235; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n22137; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n22138; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n22139; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n21920; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n22154; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n22130; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n22236; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n22237; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n22238; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n22286_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n22287_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n22288_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n22239; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n22240; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n22132; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n21970_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n21943_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n21736_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n22222; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n22223; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n22232; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n22233; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n21734_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n21735_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n22131; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n22136; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n22133; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n22134; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n22135; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n22144; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n22145; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n22140; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n22141; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n22142; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n22143; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n22224; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n22225; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n22231; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n22146; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n22147; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n22148; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n21919; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n22149; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n22150; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n22151; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n22152; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n22153; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n22290_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n22292_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n22293_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n22294_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n22296_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n22298_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n22300_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n22302_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n22304_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n22306_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n22308_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n22155; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n22156; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n22157; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n22070; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n22071; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n22072; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n22230; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n22158; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n22159; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n21913; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n21914; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n21402_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n21403_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n21442_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:191:8  */
  assign dp_wr_fork = n21443_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n21404_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n21444_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n21445_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n21446_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n21447_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n21448_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n21449_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n21450_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n21405_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n21406_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n21407_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n21408_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n21409_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n21410_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n21411_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n21412_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n21413_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n21414_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n21696_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n21415_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n21416_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n21452_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n21455_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n22309_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n22310_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n22311_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n22314_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n22315_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n22316_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n22317_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n22318_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n22319_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n22320_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n22321_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n22322_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n22323_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n22324_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n22326_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n22328_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n22330_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:238:8  */
  assign dp_wr_fork_r = n22332_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n22333_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n22334_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n22336_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n22338_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n22342_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n22344_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n22346_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n22348_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n22350_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n22352_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n22354_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n22358_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n22362_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n22364_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n22366_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n22368_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n22370_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n22372_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n22374_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n22375_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n22376_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n22377_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n21720_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n21381_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n22087; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n22088; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n22089; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n22090; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n22091; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n22092; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n22085; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n22086; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n22093; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n22094; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n22095; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n22096; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n22097; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n21259_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n21260_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n21261_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n22379_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n22380_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n22381_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n22382_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n22383_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n22384_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n22385_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n22386_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n22387_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n22388_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n22389_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n22390_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n22391_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n22392_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n22393_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n22394_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n22395_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n22397_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n22398_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n22400_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n22401_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n22402_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n22403_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n22404_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n22405_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n22406_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n22407_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n22408_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n22409_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n22410_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n22411_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n22412_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n22413_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n22414_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n22415_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n22416_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n22417_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n22418_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n22419_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n22420_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n22421_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n22422_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n22423_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n22424_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n22425_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n21259_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n21260_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n21261_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n21264_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n21352_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n21353_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n21354_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n21355_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n21358_o = n21355_o ? 3'b001 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n21360_o = n21354_o + n21352_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n21361_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n21362_o = n21361_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n21363_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n21364_o = n21363_o & n21362_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n21365_o = n21352_o & n21354_o;
  /* ../../HW/src/pcore/pcore.vhd:215:8  */
  assign n21366_o = {n21358_o, 2'b00};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n21367_o = n21352_o & n21366_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n21368_o = n21365_o == n21367_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n21369_o = n21368_o & n21353_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n21370_o = ~n21353_o;
  /* ../../HW/src/pcore/pcore.vhd:106:8  */
  assign n21371_o = {n21358_o, 2'b00};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n21372_o = $unsigned(n21371_o) >= $unsigned(n21354_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n21373_o = n21372_o & n21370_o;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n21374_o = {n21358_o, 2'b00};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n21375_o = $unsigned(n21374_o) <= $unsigned(n21360_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n21376_o = n21375_o & n21373_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n21377_o = n21369_o | n21376_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n21378_o = n21377_o & n21364_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n21381_o = n21378_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n21387_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n21389_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n21391_o = n21389_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n21393_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n21394_o = n21393_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n21395_o = dp_read_gen_valid_in_r & n21394_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n21397_o = n21395_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n21399_o = n21395_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n21401_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21402_o = n21387_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21403_o = n21387_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21404_o = n21387_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21405_o = n21387_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21406_o = n21387_o ? n21391_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21407_o = n21387_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21408_o = n21387_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21409_o = n21387_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21410_o = n21387_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21411_o = n21387_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21412_o = n21387_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21413_o = n21387_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21414_o = n21387_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21415_o = n21387_o ? n21397_o : n21401_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n21416_o = n21387_o ? n21399_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n21421_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n21422_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n21423_o = dp_write_in_r & n21422_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n21424_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n21425_o = n21423_o & n21424_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n21427_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n21429_o = n21427_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n21431_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n21432_o = n21431_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n21433_o = dp_write_gen_valid_in_r & n21432_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n21435_o = n21433_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n21439_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n21441_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21442_o = n21421_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21443_o = n21421_o ? dp_wr_fork_in_r : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21444_o = n21421_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21445_o = n21421_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21446_o = n21421_o ? n21425_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21447_o = n21421_o ? n21429_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21448_o = n21421_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21449_o = n21421_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21450_o = n21421_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21452_o = n21421_o ? n21435_o : n21439_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n21455_o = n21421_o ? 3'b000 : n21441_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n21460_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n21463_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n21464_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n21465_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n21467_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n21468_o = n21464_o ? n21465_o : n21467_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n21470_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n21471_o = n21463_o ? n21468_o : n21470_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n21473_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n21537_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n21606_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n21609_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n21610_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n21611_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n21613_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n21614_o = n21610_o ? n21611_o : n21613_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n21616_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n21617_o = n21609_o ? n21614_o : n21616_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n21619_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n21620_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n21621_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n21631_o = n21619_o ? n21620_o : n21621_o;
  assign n21673_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n21674_o = n21606_o ? 12'b000000000000 : n21673_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n21688_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n21690_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n21691_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n21692_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n21693_o = n21690_o ? n21691_o : n21692_o;
  assign n21695_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n21693_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n21696_o = n21688_o ? n21695_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n21702_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n21703_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n21704_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n21706_o = n21702_o == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n21707_o = n21706_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n21709_o = n21703_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n21710_o = n21709_o & n21707_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n21713_o = n21710_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n21715_o = n21702_o == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n21716_o = n21715_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n21719_o = n21716_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n21720_o = n21704_o ? n21713_o : n21719_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n21722_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n21724_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n21726_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n21728_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n21734_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n21735_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n21736_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n21739_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n21740_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n21742_o = n21739_o ? 96'bZ : n21740_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n21744_o = n21739_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n21749_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n21800_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n21803_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n21804_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n21805_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n21807_o = n21804_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n21808_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n21810_o = n21804_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n21811_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n21813_o = n21804_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n21814_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n21816_o = n21804_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n21817_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n21819_o = n21804_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n21820_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n21822_o = n21804_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n21823_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n21825_o = n21804_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n21826_o = dp_readdata_vm[11:0];
  assign n21827_o = {n21825_o, n21822_o, n21819_o, n21816_o, n21813_o, n21810_o, n21807_o};
  assign n21828_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21829_o = n21828_o;
      7'b0100000: n21829_o = n21828_o;
      7'b0010000: n21829_o = n21828_o;
      7'b0001000: n21829_o = n21828_o;
      7'b0000100: n21829_o = n21828_o;
      7'b0000010: n21829_o = n21828_o;
      7'b0000001: n21829_o = n21828_o;
      default: n21829_o = n21826_o;
    endcase
  assign n21830_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21831_o = n21823_o;
      7'b0100000: n21831_o = n21830_o;
      7'b0010000: n21831_o = n21830_o;
      7'b0001000: n21831_o = n21830_o;
      7'b0000100: n21831_o = n21830_o;
      7'b0000010: n21831_o = n21830_o;
      7'b0000001: n21831_o = n21830_o;
      default: n21831_o = n21830_o;
    endcase
  assign n21832_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21833_o = n21832_o;
      7'b0100000: n21833_o = n21820_o;
      7'b0010000: n21833_o = n21832_o;
      7'b0001000: n21833_o = n21832_o;
      7'b0000100: n21833_o = n21832_o;
      7'b0000010: n21833_o = n21832_o;
      7'b0000001: n21833_o = n21832_o;
      default: n21833_o = n21832_o;
    endcase
  assign n21834_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21835_o = n21834_o;
      7'b0100000: n21835_o = n21834_o;
      7'b0010000: n21835_o = n21817_o;
      7'b0001000: n21835_o = n21834_o;
      7'b0000100: n21835_o = n21834_o;
      7'b0000010: n21835_o = n21834_o;
      7'b0000001: n21835_o = n21834_o;
      default: n21835_o = n21834_o;
    endcase
  assign n21836_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21837_o = n21836_o;
      7'b0100000: n21837_o = n21836_o;
      7'b0010000: n21837_o = n21836_o;
      7'b0001000: n21837_o = n21814_o;
      7'b0000100: n21837_o = n21836_o;
      7'b0000010: n21837_o = n21836_o;
      7'b0000001: n21837_o = n21836_o;
      default: n21837_o = n21836_o;
    endcase
  assign n21838_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21839_o = n21838_o;
      7'b0100000: n21839_o = n21838_o;
      7'b0010000: n21839_o = n21838_o;
      7'b0001000: n21839_o = n21838_o;
      7'b0000100: n21839_o = n21811_o;
      7'b0000010: n21839_o = n21838_o;
      7'b0000001: n21839_o = n21838_o;
      default: n21839_o = n21838_o;
    endcase
  assign n21840_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21841_o = n21840_o;
      7'b0100000: n21841_o = n21840_o;
      7'b0010000: n21841_o = n21840_o;
      7'b0001000: n21841_o = n21840_o;
      7'b0000100: n21841_o = n21840_o;
      7'b0000010: n21841_o = n21808_o;
      7'b0000001: n21841_o = n21840_o;
      default: n21841_o = n21840_o;
    endcase
  assign n21842_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n21827_o)
      7'b1000000: n21843_o = n21842_o;
      7'b0100000: n21843_o = n21842_o;
      7'b0010000: n21843_o = n21842_o;
      7'b0001000: n21843_o = n21842_o;
      7'b0000100: n21843_o = n21842_o;
      7'b0000010: n21843_o = n21842_o;
      7'b0000001: n21843_o = n21805_o;
      default: n21843_o = n21842_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n21845_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n21848_o = n21845_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n21849_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n21850_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n21851_o = {n21843_o, n21841_o, n21839_o, n21837_o, n21835_o, n21833_o, n21831_o, n21829_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n21852_o = n21803_o ? n21851_o : n21849_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n21853_o = n21803_o ? dp_readdata2_r : n21850_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n21855_o = n21803_o ? n21848_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n21857_o = n21803_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n21859_o = n21803_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n21864_o = dp_readena_vm ? n21855_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n21913 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n21914 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n21919 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n21920 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n21927_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n21929_o = dp_rd_pid == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n21930_o = n21929_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n21932_o = dp_rd_cid == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n21933_o = n21932_o & n21930_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n21936_o = n21933_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n21938_o = dp_rd_pid == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n21939_o = n21938_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n21942_o = n21939_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n21943_o = n21927_o ? n21936_o : n21942_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n21951_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n21952_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n21953_o = dp_mcast_addr + n21951_o;
  /* ../../HW/src/pcore/pcore.vhd:1022:1  */
  assign n21956_o = dp_wr_fork ? 5'b00000 : 5'b00100;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n21957_o = n21951_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n21958_o = n21951_o & n21956_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n21959_o = n21957_o == n21958_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n21960_o = n21959_o & n21952_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n21961_o = ~n21952_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n21962_o = $unsigned(n21956_o) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n21963_o = n21962_o & n21961_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n21964_o = $unsigned(n21956_o) <= $unsigned(n21953_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n21965_o = n21964_o & n21963_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n21966_o = n21960_o | n21965_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n21967_o = n21966_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n21970_o = n21967_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n21972_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n21973_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n21974_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n21975 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n21976 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n21977 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n21972_o),
    .x1_in(n21973_o),
    .x2_in(n21974_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n21984_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n21985_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n21986_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n21987 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n21988 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n21989 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n21984_o),
    .x1_in(n21985_o),
    .x2_in(n21986_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n21996_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n21997_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n21998_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n21999 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n22000 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n22001 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n21996_o),
    .x1_in(n21997_o),
    .x2_in(n21998_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n22008_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n22009_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n22010_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n22011 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n22012 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n22013 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n22008_o),
    .x1_in(n22009_o),
    .x2_in(n22010_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n22020_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n22021_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n22022_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n22023 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n22024 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n22025 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n22020_o),
    .x1_in(n22021_o),
    .x2_in(n22022_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n22032_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n22033_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n22034_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n22035 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n22036 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n22037 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n22032_o),
    .x1_in(n22033_o),
    .x2_in(n22034_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n22044_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n22045_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n22046_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n22047 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n22048 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n22049 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n22044_o),
    .x1_in(n22045_o),
    .x2_in(n22046_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n22056_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n22057_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n22058_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n22059 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n22060 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n22061 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n22056_o),
    .x1_in(n22057_o),
    .x2_in(n22058_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n22068_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n22069_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n22070 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n22071 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n22072 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n22081 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n22082 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n22083_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n22084_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n22085 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n22086 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n22087 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n22088 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n22089 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n22090 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n22091 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n22092 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n22093 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n22094 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n22095 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n22096 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n22097 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n22083_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n22084_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n22130 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n22131 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n22132 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n22133 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n22134 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n22135 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n22136 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n22137 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n22138 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n22139 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n22140 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n22141 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n22142 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n22143 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n22144 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n22145 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n22146 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n22147 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n22148 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n22149 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n22150 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n22151 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n22152 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n22153 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n22154 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n22155 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n22156 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n22157 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n22158 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n22159 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_1_0 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n22220 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n22221 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n22222 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n22223 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n22224 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n22225 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n22226 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n22227 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n22228 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n22229 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n22230 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n22231 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n22232 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n22233 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n22234 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n22235 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n22236 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n22237 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n22238 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n22239 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n22240 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n22286_o = {alu_7_i_n22059, alu_6_i_n22047, alu_5_i_n22035, alu_4_i_n22023, alu_3_i_n22011, alu_2_i_n21999, alu_1_i_n21987, alu_0_i_n21975};
  assign n22287_o = {alu_7_i_n22061, alu_6_i_n22049, alu_5_i_n22037, alu_4_i_n22025, alu_3_i_n22013, alu_2_i_n22001, alu_1_i_n21989, alu_0_i_n21977};
  assign n22288_o = {alu_7_i_n22060, alu_6_i_n22048, alu_5_i_n22036, alu_4_i_n22024, alu_3_i_n22012, alu_2_i_n22000, alu_1_i_n21988, alu_0_i_n21976};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22289_o = dp_readena_vm ? n21852_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22290_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n22290_q <= n22289_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22291_o = dp_readena_vm ? n21853_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22292_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n22292_q <= n22291_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22293_q <= 1'b0;
    else
      n22293_q <= n21864_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22294_q <= 1'b0;
    else
      n22294_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22295_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22296_q <= 1'b0;
    else
      n22296_q <= n22295_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22297_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22298_q <= 2'b00;
    else
      n22298_q <= n22297_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22299_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22300_q <= 2'b00;
    else
      n22300_q <= n22299_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22301_o = dp_readena_vm ? n21857_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22302_q <= 3'b000;
    else
      n22302_q <= n22301_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22303_o = dp_readena_vm ? n21859_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22304_q <= 3'b000;
    else
      n22304_q <= n22303_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22305_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22306_q <= 1'b0;
    else
      n22306_q <= n22305_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n22307_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n21800_o)
    if (n21800_o)
      n22308_q <= 2'b00;
    else
      n22308_q <= n22307_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22309_q <= 3'b000;
    else
      n22309_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22310_q <= 3'b000;
    else
      n22310_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22311_q <= 2'b00;
    else
      n22311_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22314_q <= 3'b000;
    else
      n22314_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22315_q <= 3'b000;
    else
      n22315_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22316_q <= 1'b0;
    else
      n22316_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22317_q <= 2'b00;
    else
      n22317_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22318_q <= 2'b00;
    else
      n22318_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22319_q <= 1'b0;
    else
      n22319_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22320_q <= 2'b00;
    else
      n22320_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22321_q <= 22'b0000000000000000000000;
    else
      n22321_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22322_q <= 3'b000;
    else
      n22322_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22323_q <= 22'b0000000000000000000000;
    else
      n22323_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22324_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n22324_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22325_o = n21473_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22326_q <= 1'b0;
    else
      n22326_q <= n22325_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22327_o = n21473_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22328_q <= 1'b0;
    else
      n22328_q <= n22327_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22329_o = n21619_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22330_q <= 1'b0;
    else
      n22330_q <= n22329_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22331_o = n21619_o ? dp_wr_fork : dp_wr_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22332_q <= 1'b0;
    else
      n22332_q <= n22331_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22333_q <= 22'b0000000000000000000000;
    else
      n22333_q <= n21471_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22334_q <= 22'b0000000000000000000000;
    else
      n22334_q <= n21617_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22335_o = n21619_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22336_q <= 6'b000000;
    else
      n22336_q <= n22335_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22337_o = n21619_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22338_q <= 1'b0;
    else
      n22338_q <= n22337_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22341_o = n21619_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22342_q <= 3'b000;
    else
      n22342_q <= n22341_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22343_o = n21619_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22344_q <= 2'b00;
    else
      n22344_q <= n22343_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22345_o = n21619_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22346_q <= 1'b0;
    else
      n22346_q <= n22345_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n22347_o = n21619_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22348_q <= 22'b0000000000000000000000;
    else
      n22348_q <= n22347_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22349_o = n21473_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22350_q <= 1'b0;
    else
      n22350_q <= n22349_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22351_o = n21473_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22352_q <= 3'b000;
    else
      n22352_q <= n22351_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22353_o = n21473_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22354_q <= 2'b00;
    else
      n22354_q <= n22353_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n22355_o = ~n21460_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n22356_o = n21473_o & n22355_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22357_o = n22356_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n22358_q <= n22357_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n22359_o = ~n21460_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n22360_o = n21473_o & n22359_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22361_o = n22360_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n22362_q <= n22361_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22363_o = n21473_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22364_q <= 1'b0;
    else
      n22364_q <= n22363_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22365_o = n21473_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22366_q <= 2'b00;
    else
      n22366_q <= n22365_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22367_o = n21473_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22368_q <= 2'b00;
    else
      n22368_q <= n22367_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22369_o = n21473_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22370_q <= 1'b0;
    else
      n22370_q <= n22369_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n22371_o = n21473_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22372_q <= 2'b00;
    else
      n22372_q <= n22371_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22373_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n22373_q <= n21631_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n22374_o = {n21674_o, n22373_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22375_q <= 3'b000;
    else
      n22375_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n21460_o)
    if (n21460_o)
      n22376_q <= 3'b000;
    else
      n22376_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n21606_o)
    if (n21606_o)
      n22377_q <= 3'b000;
    else
      n22377_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22379_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n22379_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22380_q <= 32'b00000000000000000000000000000000;
    else
      n22380_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22381_q <= 1'b0;
    else
      n22381_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22382_q <= 1'b0;
    else
      n22382_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22383_q <= 1'b0;
    else
      n22383_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22384_q <= 2'b00;
    else
      n22384_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22385_q <= 4'b0000;
    else
      n22385_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22386_q <= 1'b0;
    else
      n22386_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22387_q <= 4'b0000;
    else
      n22387_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22388_q <= 1'b0;
    else
      n22388_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22389_q <= 4'b0000;
    else
      n22389_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22390_q <= 1'b0;
    else
      n22390_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22391_q <= 1'b0;
    else
      n22391_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22392_q <= 2'b00;
    else
      n22392_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n21749_o)
    if (n21749_o)
      n22393_q <= 28'b0000000000000000000000000000;
    else
      n22393_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22394_q <= 1'b0;
    else
      n22394_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22395_q <= 1'b0;
    else
      n22395_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22397_q <= 1'b0;
    else
      n22397_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n21537_o)
    if (n21537_o)
      n22398_q <= 1'b0;
    else
      n22398_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22400_q <= 1'b0;
    else
      n22400_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22401_q <= 1'b0;
    else
      n22401_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22402_q <= 1'b0;
    else
      n22402_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22403_q <= 22'b0000000000000000000000;
    else
      n22403_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22404_q <= 1'b0;
    else
      n22404_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22405_q <= 22'b0000000000000000000000;
    else
      n22405_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22406_q <= 22'b0000000000000000000000;
    else
      n22406_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22407_q <= 1'b0;
    else
      n22407_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22408_q <= 22'b0000000000000000000000;
    else
      n22408_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22409_q <= 6'b000000;
    else
      n22409_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22410_q <= 1'b0;
    else
      n22410_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22411_q <= 1'b0;
    else
      n22411_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22412_q <= 1'b0;
    else
      n22412_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22413_q <= 3'b000;
    else
      n22413_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22414_q <= 2'b00;
    else
      n22414_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22415_q <= 1'b0;
    else
      n22415_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22416_q <= 1'b0;
    else
      n22416_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22417_q <= 3'b000;
    else
      n22417_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22418_q <= 2'b00;
    else
      n22418_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22419_q <= 1'b0;
    else
      n22419_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22420_q <= 2'b00;
    else
      n22420_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22421_q <= 2'b00;
    else
      n22421_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22422_q <= 1'b0;
    else
      n22422_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22423_q <= 2'b00;
    else
      n22423_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22424_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n22424_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n21264_o)
    if (n21264_o)
      n22425_q <= 1'b0;
    else
      n22425_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n22426_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n22427_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_0_3
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n20077_o;
  wire n20078_o;
  wire n20079_o;
  wire n20082_o;
  wire [4:0] n20170_o;
  wire n20171_o;
  wire [4:0] n20172_o;
  wire n20173_o;
  wire [2:0] n20176_o;
  wire [4:0] n20178_o;
  wire n20179_o;
  wire n20180_o;
  wire n20181_o;
  wire n20182_o;
  wire [4:0] n20183_o;
  wire [4:0] n20184_o;
  wire [4:0] n20185_o;
  wire n20186_o;
  wire n20187_o;
  wire n20188_o;
  wire [4:0] n20189_o;
  wire n20190_o;
  wire n20191_o;
  wire [4:0] n20192_o;
  wire n20193_o;
  wire n20194_o;
  wire n20195_o;
  wire n20196_o;
  wire n20199_o;
  wire n20205_o;
  wire n20207_o;
  wire [2:0] n20209_o;
  wire n20211_o;
  wire n20212_o;
  wire n20213_o;
  wire [2:0] n20215_o;
  wire [2:0] n20217_o;
  wire [2:0] n20219_o;
  wire n20220_o;
  wire n20221_o;
  wire [21:0] n20222_o;
  wire n20223_o;
  wire [2:0] n20224_o;
  wire [1:0] n20225_o;
  wire n20226_o;
  wire [21:0] n20227_o;
  wire n20228_o;
  wire [1:0] n20229_o;
  wire [1:0] n20230_o;
  wire n20231_o;
  wire [1:0] n20232_o;
  wire [2:0] n20233_o;
  wire [2:0] n20234_o;
  wire n20239_o;
  wire n20240_o;
  wire n20241_o;
  wire n20242_o;
  wire n20243_o;
  wire n20245_o;
  wire [2:0] n20247_o;
  wire n20249_o;
  wire n20250_o;
  wire n20251_o;
  wire [2:0] n20253_o;
  wire [2:0] n20257_o;
  wire [2:0] n20259_o;
  wire n20260_o;
  wire [21:0] n20262_o;
  wire [5:0] n20263_o;
  wire n20264_o;
  wire [2:0] n20265_o;
  wire [1:0] n20266_o;
  wire n20267_o;
  wire [21:0] n20268_o;
  wire [2:0] n20270_o;
  wire [2:0] n20273_o;
  wire n20278_o;
  wire n20281_o;
  wire n20282_o;
  wire [21:0] n20283_o;
  wire [21:0] n20285_o;
  wire [21:0] n20286_o;
  wire [21:0] n20288_o;
  wire [21:0] n20289_o;
  wire n20291_o;
  wire n20355_o;
  wire n20424_o;
  wire n20427_o;
  wire n20428_o;
  wire [21:0] n20429_o;
  wire [21:0] n20431_o;
  wire [21:0] n20432_o;
  wire [21:0] n20434_o;
  wire [21:0] n20435_o;
  wire n20437_o;
  wire [83:0] n20438_o;
  wire [83:0] n20439_o;
  wire [83:0] n20449_o;
  wire [11:0] n20491_o;
  wire [11:0] n20492_o;
  wire n20506_o;
  wire n20508_o;
  wire [11:0] n20509_o;
  wire [11:0] n20510_o;
  wire [11:0] n20511_o;
  wire [95:0] n20513_o;
  wire [95:0] n20514_o;
  wire [1:0] n20520_o;
  wire [2:0] n20521_o;
  wire n20522_o;
  wire n20524_o;
  wire n20525_o;
  wire n20527_o;
  wire n20528_o;
  wire n20531_o;
  wire n20533_o;
  wire n20534_o;
  wire n20537_o;
  wire n20538_o;
  wire [1:0] n20540_o;
  wire [1:0] n20542_o;
  wire n20544_o;
  wire [1:0] n20546_o;
  wire [1:0] n20552_o;
  wire [2:0] n20553_o;
  wire [4:0] n20554_o;
  wire n20557_o;
  wire [95:0] n20558_o;
  wire [95:0] n20560_o;
  wire n20562_o;
  wire n20567_o;
  wire n20618_o;
  wire n20621_o;
  wire [2:0] n20622_o;
  wire [11:0] n20623_o;
  wire n20625_o;
  wire [11:0] n20626_o;
  wire n20628_o;
  wire [11:0] n20629_o;
  wire n20631_o;
  wire [11:0] n20632_o;
  wire n20634_o;
  wire [11:0] n20635_o;
  wire n20637_o;
  wire [11:0] n20638_o;
  wire n20640_o;
  wire [11:0] n20641_o;
  wire n20643_o;
  wire [11:0] n20644_o;
  wire [6:0] n20645_o;
  wire [11:0] n20646_o;
  reg [11:0] n20647_o;
  wire [11:0] n20648_o;
  reg [11:0] n20649_o;
  wire [11:0] n20650_o;
  reg [11:0] n20651_o;
  wire [11:0] n20652_o;
  reg [11:0] n20653_o;
  wire [11:0] n20654_o;
  reg [11:0] n20655_o;
  wire [11:0] n20656_o;
  reg [11:0] n20657_o;
  wire [11:0] n20658_o;
  reg [11:0] n20659_o;
  wire [11:0] n20660_o;
  reg [11:0] n20661_o;
  wire n20663_o;
  wire n20666_o;
  wire [95:0] n20667_o;
  wire [95:0] n20668_o;
  wire [95:0] n20669_o;
  wire [95:0] n20670_o;
  wire [95:0] n20671_o;
  wire n20673_o;
  wire [2:0] n20675_o;
  wire [2:0] n20677_o;
  wire n20682_o;
  wire [12:0] xregister_file_i_n20731;
  wire [255:0] xregister_file_i_n20732;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n20737;
  wire [12:0] iregister_i_n20738;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n20745_o;
  wire n20747_o;
  wire n20748_o;
  wire n20750_o;
  wire n20751_o;
  wire n20754_o;
  wire n20756_o;
  wire n20757_o;
  wire n20760_o;
  wire n20761_o;
  wire [4:0] n20769_o;
  wire n20770_o;
  wire [4:0] n20771_o;
  wire [4:0] n20772_o;
  wire [4:0] n20774_o;
  wire n20775_o;
  wire n20776_o;
  wire n20777_o;
  wire n20779_o;
  wire n20780_o;
  wire n20782_o;
  wire n20783_o;
  wire n20784_o;
  wire n20785_o;
  wire n20788_o;
  wire [31:0] n20791_o;
  wire [11:0] n20792_o;
  wire [11:0] n20793_o;
  wire [31:0] alu_0_i_n20794;
  wire alu_0_i_n20795;
  wire [11:0] alu_0_i_n20796;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n20803_o;
  wire [11:0] n20804_o;
  wire [11:0] n20805_o;
  wire [31:0] alu_1_i_n20806;
  wire alu_1_i_n20807;
  wire [11:0] alu_1_i_n20808;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n20815_o;
  wire [11:0] n20816_o;
  wire [11:0] n20817_o;
  wire [31:0] alu_2_i_n20818;
  wire alu_2_i_n20819;
  wire [11:0] alu_2_i_n20820;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n20827_o;
  wire [11:0] n20828_o;
  wire [11:0] n20829_o;
  wire [31:0] alu_3_i_n20830;
  wire alu_3_i_n20831;
  wire [11:0] alu_3_i_n20832;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n20839_o;
  wire [11:0] n20840_o;
  wire [11:0] n20841_o;
  wire [31:0] alu_4_i_n20842;
  wire alu_4_i_n20843;
  wire [11:0] alu_4_i_n20844;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n20851_o;
  wire [11:0] n20852_o;
  wire [11:0] n20853_o;
  wire [31:0] alu_5_i_n20854;
  wire alu_5_i_n20855;
  wire [11:0] alu_5_i_n20856;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n20863_o;
  wire [11:0] n20864_o;
  wire [11:0] n20865_o;
  wire [31:0] alu_6_i_n20866;
  wire alu_6_i_n20867;
  wire [11:0] alu_6_i_n20868;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n20875_o;
  wire [11:0] n20876_o;
  wire [11:0] n20877_o;
  wire [31:0] alu_7_i_n20878;
  wire alu_7_i_n20879;
  wire [11:0] alu_7_i_n20880;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n20887_o;
  wire n20888_o;
  wire [12:0] ialu_i_n20889;
  wire ialu_i_n20890;
  wire ialu_i_n20891;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n20900;
  wire [95:0] register_bank_i_n20901;
  wire [16:0] n20902_o;
  wire [16:0] n20903_o;
  wire [95:0] register_bank_i_n20904;
  wire register_bank_i_n20905;
  wire register_bank_i_n20906;
  wire [2:0] register_bank_i_n20907;
  wire [2:0] register_bank_i_n20908;
  wire [1:0] register_bank_i_n20909;
  wire [2:0] register_bank_i_n20910;
  wire [2:0] register_bank_i_n20911;
  wire register_bank_i_n20912;
  wire [1:0] register_bank_i_n20913;
  wire [1:0] register_bank_i_n20914;
  wire register_bank_i_n20915;
  wire [1:0] register_bank_i_n20916;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n20949;
  wire instr_decoder2_i_n20950;
  wire [3:0] instr_decoder2_i_n20951;
  wire instr_decoder2_i_n20952;
  wire instr_decoder2_i_n20953;
  wire instr_decoder2_i_n20954;
  wire instr_decoder2_i_n20955;
  wire [11:0] instr_decoder2_i_n20956;
  wire [11:0] instr_decoder2_i_n20957;
  wire [11:0] instr_decoder2_i_n20958;
  wire instr_decoder2_i_n20959;
  wire instr_decoder2_i_n20960;
  wire instr_decoder2_i_n20961;
  wire [7:0] instr_decoder2_i_n20962;
  wire instr_decoder2_i_n20963;
  wire [11:0] instr_decoder2_i_n20964;
  wire instr_decoder2_i_n20965;
  wire instr_decoder2_i_n20966;
  wire [3:0] instr_decoder2_i_n20967;
  wire [3:0] instr_decoder2_i_n20968;
  wire instr_decoder2_i_n20969;
  wire instr_decoder2_i_n20970;
  wire [2:0] instr_decoder2_i_n20971;
  wire [12:0] instr_decoder2_i_n20972;
  wire instr_decoder2_i_n20973;
  wire [4:0] instr_decoder2_i_n20974;
  wire [12:0] instr_decoder2_i_n20975;
  wire [12:0] instr_decoder2_i_n20976;
  wire [7:0] instr_decoder2_i_n20977;
  wire [7:0] instr_decoder2_i_n20978;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n21039;
  wire instr_dispatch2_i1_n21040;
  wire [11:0] instr_dispatch2_i1_n21041;
  wire [11:0] instr_dispatch2_i1_n21042;
  wire instr_dispatch2_i1_n21043;
  wire instr_dispatch2_i1_n21044;
  wire instr_dispatch2_i1_n21045;
  wire instr_dispatch2_i1_n21046;
  wire instr_dispatch2_i1_n21047;
  wire instr_dispatch2_i1_n21048;
  wire instr_dispatch2_i1_n21049;
  wire instr_dispatch2_i1_n21050;
  wire [11:0] instr_dispatch2_i1_n21051;
  wire [7:0] instr_dispatch2_i1_n21052;
  wire [95:0] instr_dispatch2_i1_n21053;
  wire [7:0] instr_dispatch2_i1_n21054;
  wire [95:0] instr_dispatch2_i1_n21055;
  wire [95:0] instr_dispatch2_i1_n21056;
  wire [11:0] instr_dispatch2_i1_n21057;
  wire [4:0] instr_dispatch2_i1_n21058;
  wire [3:0] instr_dispatch2_i1_n21059;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n21105_o;
  wire [95:0] n21106_o;
  wire [7:0] n21107_o;
  wire [95:0] n21108_o;
  reg [95:0] n21109_q;
  wire [95:0] n21110_o;
  reg [95:0] n21111_q;
  reg n21112_q;
  reg n21113_q;
  wire n21114_o;
  reg n21115_q;
  wire [1:0] n21116_o;
  reg [1:0] n21117_q;
  wire [1:0] n21118_o;
  reg [1:0] n21119_q;
  wire [2:0] n21120_o;
  reg [2:0] n21121_q;
  wire [2:0] n21122_o;
  reg [2:0] n21123_q;
  wire n21124_o;
  reg n21125_q;
  wire [1:0] n21126_o;
  reg [1:0] n21127_q;
  reg [2:0] n21128_q;
  reg [2:0] n21129_q;
  reg [1:0] n21130_q;
  reg [2:0] n21133_q;
  reg [2:0] n21134_q;
  reg n21135_q;
  reg [1:0] n21136_q;
  reg [1:0] n21137_q;
  reg n21138_q;
  reg [1:0] n21139_q;
  reg [21:0] n21140_q;
  reg [2:0] n21141_q;
  reg [21:0] n21142_q;
  reg [95:0] n21143_q;
  wire n21144_o;
  reg n21145_q;
  wire n21146_o;
  reg n21147_q;
  wire n21148_o;
  reg n21149_q;
  reg [21:0] n21152_q;
  reg [21:0] n21153_q;
  wire [5:0] n21154_o;
  reg [5:0] n21155_q;
  wire n21156_o;
  reg n21157_q;
  wire [2:0] n21160_o;
  reg [2:0] n21161_q;
  wire [1:0] n21162_o;
  reg [1:0] n21163_q;
  wire n21164_o;
  reg n21165_q;
  wire [21:0] n21166_o;
  reg [21:0] n21167_q;
  wire n21168_o;
  reg n21169_q;
  wire [2:0] n21170_o;
  reg [2:0] n21171_q;
  wire [1:0] n21172_o;
  reg [1:0] n21173_q;
  wire n21174_o;
  wire n21175_o;
  wire n21176_o;
  reg n21177_q;
  wire n21178_o;
  wire n21179_o;
  wire [21:0] n21180_o;
  reg [21:0] n21181_q;
  wire n21182_o;
  reg n21183_q;
  wire [1:0] n21184_o;
  reg [1:0] n21185_q;
  wire [1:0] n21186_o;
  reg [1:0] n21187_q;
  wire n21188_o;
  reg n21189_q;
  wire [1:0] n21190_o;
  reg [1:0] n21191_q;
  reg [83:0] n21192_q;
  wire [95:0] n21193_o;
  reg [2:0] n21194_q;
  reg [2:0] n21195_q;
  reg [2:0] n21196_q;
  reg [79:0] n21198_q;
  reg [31:0] n21199_q;
  reg n21200_q;
  reg n21201_q;
  reg n21202_q;
  reg [1:0] n21203_q;
  reg [3:0] n21204_q;
  reg n21205_q;
  reg [3:0] n21206_q;
  reg n21207_q;
  reg [3:0] n21208_q;
  reg n21209_q;
  reg n21210_q;
  reg [1:0] n21211_q;
  reg [27:0] n21212_q;
  reg n21213_q;
  reg n21214_q;
  reg n21216_q;
  reg n21217_q;
  reg n21219_q;
  reg n21220_q;
  reg n21221_q;
  reg [21:0] n21222_q;
  reg n21223_q;
  reg [21:0] n21224_q;
  reg [21:0] n21225_q;
  reg n21226_q;
  reg [21:0] n21227_q;
  reg [5:0] n21228_q;
  reg n21229_q;
  reg n21230_q;
  reg n21231_q;
  reg [2:0] n21232_q;
  reg [1:0] n21233_q;
  reg n21234_q;
  reg n21235_q;
  reg [2:0] n21236_q;
  reg [1:0] n21237_q;
  reg n21238_q;
  reg [1:0] n21239_q;
  reg [1:0] n21240_q;
  reg n21241_q;
  reg [1:0] n21242_q;
  reg [95:0] n21243_q;
  reg n21244_q;
  wire [2:0] n21245_o;
  wire [2:0] n21246_o;
  assign i_y_neg_out = n20887_o;
  assign i_y_zero_out = n20888_o;
  assign dp_readdata_out = n20560_o;
  assign dp_readdata_vm_out = n20562_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n21245_o;
  assign dp_read_vaddr_out = n21246_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n20540_o;
  assign dp_read_data_type_out = n20542_o;
  assign dp_read_stream_out = n20544_o;
  assign dp_read_stream_id_out = n20546_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n20900; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n20901; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n21039; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n21040; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n21048; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n21045; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n21046; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n21047; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n21053; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n21054; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n20956; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n20957; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n20958; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n20738; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n20973; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n20949; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n21055; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n21056; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n21057; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n21105_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n21106_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n21107_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n21058; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n21059; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n20951; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n20788_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n20761_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n20554_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n21041; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n21042; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n21051; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n21052; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n20552_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n20553_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n20950; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n20955; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n20952; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n20953; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n20954; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n20963; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n20964; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n20959; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n20960; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n20961; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n20962; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n21043; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n21044; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n21050; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n20965; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n20966; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n20967; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n20737; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n20968; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n20969; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n20970; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n20971; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n20972; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n21109_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n21111_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n21112_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n21113_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n21115_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n21117_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n21119_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n21121_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n21123_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n21125_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n21127_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n20974; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n20975; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n20976; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n20889; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n20890; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n20891; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n21049; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n20977; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n20978; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n20731; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n20732; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n20220_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n20221_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n20260_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n20222_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n20262_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n20263_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n20264_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n20265_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n20266_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n20267_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n20268_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n20223_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n20224_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n20225_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n20226_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n20227_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n20228_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n20229_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n20230_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n20231_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n20232_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n20514_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n20233_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n20234_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n20270_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n20273_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n21128_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n21129_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n21130_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n21133_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n21134_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n21135_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n21136_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n21137_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n21138_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n21139_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n21140_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n21141_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n21142_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n21143_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n21145_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n21147_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n21149_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n21152_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n21153_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n21155_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n21157_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n21161_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n21163_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n21165_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n21167_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n21169_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n21171_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n21173_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n21177_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n21181_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n21183_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n21185_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n21187_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n21189_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n21191_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n21193_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n21194_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n21195_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n21196_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n20538_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n20199_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n20906; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n20907; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n20908; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n20909; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n20910; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n20911; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n20904; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n20905; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n20912; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n20913; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n20914; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n20915; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n20916; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n20077_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n20078_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n20079_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n21198_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n21199_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n21200_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n21201_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n21202_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n21203_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n21204_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n21205_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n21206_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n21207_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n21208_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n21209_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n21210_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n21211_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n21212_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n21213_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n21214_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n21216_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n21217_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n21219_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n21220_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n21221_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n21222_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n21223_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n21224_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n21225_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n21226_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n21227_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n21228_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n21229_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n21230_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n21231_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n21232_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n21233_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n21234_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n21235_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n21236_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n21237_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n21238_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n21239_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n21240_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n21241_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n21242_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n21243_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n21244_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n20077_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n20078_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n20079_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n20082_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n20170_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n20171_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n20172_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n20173_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n20176_o = n20173_o ? 3'b000 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n20178_o = n20172_o + n20170_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n20179_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n20180_o = n20179_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n20181_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n20182_o = n20181_o & n20180_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n20183_o = n20170_o & n20172_o;
  /* ../../HW/src/pcore/pcore.vhd:215:8  */
  assign n20184_o = {n20176_o, 2'b11};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n20185_o = n20170_o & n20184_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n20186_o = n20183_o == n20185_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n20187_o = n20186_o & n20171_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n20188_o = ~n20171_o;
  /* ../../HW/src/pcore/pcore.vhd:106:8  */
  assign n20189_o = {n20176_o, 2'b11};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n20190_o = $unsigned(n20189_o) >= $unsigned(n20172_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n20191_o = n20190_o & n20188_o;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n20192_o = {n20176_o, 2'b11};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n20193_o = $unsigned(n20192_o) <= $unsigned(n20178_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n20194_o = n20193_o & n20191_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n20195_o = n20187_o | n20194_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n20196_o = n20195_o & n20182_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n20199_o = n20196_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n20205_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n20207_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n20209_o = n20207_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n20211_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n20212_o = n20211_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n20213_o = dp_read_gen_valid_in_r & n20212_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n20215_o = n20213_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n20217_o = n20213_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n20219_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20220_o = n20205_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20221_o = n20205_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20222_o = n20205_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20223_o = n20205_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20224_o = n20205_o ? n20209_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20225_o = n20205_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20226_o = n20205_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20227_o = n20205_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20228_o = n20205_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20229_o = n20205_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20230_o = n20205_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20231_o = n20205_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20232_o = n20205_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20233_o = n20205_o ? n20215_o : n20219_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n20234_o = n20205_o ? n20217_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n20239_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n20240_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n20241_o = dp_write_in_r & n20240_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n20242_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n20243_o = n20241_o & n20242_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n20245_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n20247_o = n20245_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n20249_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n20250_o = n20249_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n20251_o = dp_write_gen_valid_in_r & n20250_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n20253_o = n20251_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n20257_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n20259_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20260_o = n20239_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20262_o = n20239_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20263_o = n20239_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20264_o = n20239_o ? n20243_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20265_o = n20239_o ? n20247_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20266_o = n20239_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20267_o = n20239_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20268_o = n20239_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20270_o = n20239_o ? n20253_o : n20257_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n20273_o = n20239_o ? 3'b000 : n20259_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n20278_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n20281_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n20282_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n20283_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n20285_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n20286_o = n20282_o ? n20283_o : n20285_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n20288_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n20289_o = n20281_o ? n20286_o : n20288_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n20291_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n20355_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n20424_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n20427_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n20428_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n20429_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n20431_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n20432_o = n20428_o ? n20429_o : n20431_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n20434_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n20435_o = n20427_o ? n20432_o : n20434_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n20437_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n20438_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n20439_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n20449_o = n20437_o ? n20438_o : n20439_o;
  assign n20491_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n20492_o = n20424_o ? 12'b000000000000 : n20491_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n20506_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n20508_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n20509_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n20510_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n20511_o = n20508_o ? n20509_o : n20510_o;
  assign n20513_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n20511_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n20514_o = n20506_o ? n20513_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n20520_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n20521_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n20522_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n20524_o = n20520_o == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n20525_o = n20524_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n20527_o = n20521_o == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n20528_o = n20527_o & n20525_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n20531_o = n20528_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n20533_o = n20520_o == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n20534_o = n20533_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n20537_o = n20534_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n20538_o = n20522_o ? n20531_o : n20537_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n20540_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n20542_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n20544_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n20546_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n20552_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n20553_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n20554_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n20557_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n20558_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n20560_o = n20557_o ? 96'bZ : n20558_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n20562_o = n20557_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n20567_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n20618_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n20621_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n20622_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n20623_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n20625_o = n20622_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n20626_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n20628_o = n20622_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n20629_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n20631_o = n20622_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n20632_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n20634_o = n20622_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n20635_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n20637_o = n20622_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n20638_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n20640_o = n20622_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n20641_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n20643_o = n20622_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n20644_o = dp_readdata_vm[11:0];
  assign n20645_o = {n20643_o, n20640_o, n20637_o, n20634_o, n20631_o, n20628_o, n20625_o};
  assign n20646_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20647_o = n20646_o;
      7'b0100000: n20647_o = n20646_o;
      7'b0010000: n20647_o = n20646_o;
      7'b0001000: n20647_o = n20646_o;
      7'b0000100: n20647_o = n20646_o;
      7'b0000010: n20647_o = n20646_o;
      7'b0000001: n20647_o = n20646_o;
      default: n20647_o = n20644_o;
    endcase
  assign n20648_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20649_o = n20641_o;
      7'b0100000: n20649_o = n20648_o;
      7'b0010000: n20649_o = n20648_o;
      7'b0001000: n20649_o = n20648_o;
      7'b0000100: n20649_o = n20648_o;
      7'b0000010: n20649_o = n20648_o;
      7'b0000001: n20649_o = n20648_o;
      default: n20649_o = n20648_o;
    endcase
  assign n20650_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20651_o = n20650_o;
      7'b0100000: n20651_o = n20638_o;
      7'b0010000: n20651_o = n20650_o;
      7'b0001000: n20651_o = n20650_o;
      7'b0000100: n20651_o = n20650_o;
      7'b0000010: n20651_o = n20650_o;
      7'b0000001: n20651_o = n20650_o;
      default: n20651_o = n20650_o;
    endcase
  assign n20652_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20653_o = n20652_o;
      7'b0100000: n20653_o = n20652_o;
      7'b0010000: n20653_o = n20635_o;
      7'b0001000: n20653_o = n20652_o;
      7'b0000100: n20653_o = n20652_o;
      7'b0000010: n20653_o = n20652_o;
      7'b0000001: n20653_o = n20652_o;
      default: n20653_o = n20652_o;
    endcase
  assign n20654_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20655_o = n20654_o;
      7'b0100000: n20655_o = n20654_o;
      7'b0010000: n20655_o = n20654_o;
      7'b0001000: n20655_o = n20632_o;
      7'b0000100: n20655_o = n20654_o;
      7'b0000010: n20655_o = n20654_o;
      7'b0000001: n20655_o = n20654_o;
      default: n20655_o = n20654_o;
    endcase
  assign n20656_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20657_o = n20656_o;
      7'b0100000: n20657_o = n20656_o;
      7'b0010000: n20657_o = n20656_o;
      7'b0001000: n20657_o = n20656_o;
      7'b0000100: n20657_o = n20629_o;
      7'b0000010: n20657_o = n20656_o;
      7'b0000001: n20657_o = n20656_o;
      default: n20657_o = n20656_o;
    endcase
  assign n20658_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20659_o = n20658_o;
      7'b0100000: n20659_o = n20658_o;
      7'b0010000: n20659_o = n20658_o;
      7'b0001000: n20659_o = n20658_o;
      7'b0000100: n20659_o = n20658_o;
      7'b0000010: n20659_o = n20626_o;
      7'b0000001: n20659_o = n20658_o;
      default: n20659_o = n20658_o;
    endcase
  assign n20660_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n20645_o)
      7'b1000000: n20661_o = n20660_o;
      7'b0100000: n20661_o = n20660_o;
      7'b0010000: n20661_o = n20660_o;
      7'b0001000: n20661_o = n20660_o;
      7'b0000100: n20661_o = n20660_o;
      7'b0000010: n20661_o = n20660_o;
      7'b0000001: n20661_o = n20623_o;
      default: n20661_o = n20660_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n20663_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n20666_o = n20663_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n20667_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n20668_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n20669_o = {n20661_o, n20659_o, n20657_o, n20655_o, n20653_o, n20651_o, n20649_o, n20647_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n20670_o = n20621_o ? n20669_o : n20667_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n20671_o = n20621_o ? dp_readdata2_r : n20668_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n20673_o = n20621_o ? n20666_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n20675_o = n20621_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n20677_o = n20621_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n20682_o = dp_readena_vm ? n20673_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n20731 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n20732 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n20737 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n20738 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n20745_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n20747_o = dp_rd_pid == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n20748_o = n20747_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n20750_o = dp_rd_cid == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n20751_o = n20750_o & n20748_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n20754_o = n20751_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n20756_o = dp_rd_pid == 2'b11;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n20757_o = n20756_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n20760_o = n20757_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n20761_o = n20745_o ? n20754_o : n20760_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n20769_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n20770_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n20771_o = dp_mcast_addr + n20769_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n20772_o = n20769_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n20774_o = n20769_o & 5'b00011;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n20775_o = n20772_o == n20774_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n20776_o = n20775_o & n20770_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n20777_o = ~n20770_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n20779_o = $unsigned(5'b00011) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n20780_o = n20779_o & n20777_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n20782_o = $unsigned(5'b00011) <= $unsigned(n20771_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n20783_o = n20782_o & n20780_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n20784_o = n20776_o | n20783_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n20785_o = n20784_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n20788_o = n20785_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n20791_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n20792_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n20793_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n20794 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n20795 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n20796 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20791_o),
    .x1_in(n20792_o),
    .x2_in(n20793_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n20803_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n20804_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n20805_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n20806 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n20807 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n20808 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20803_o),
    .x1_in(n20804_o),
    .x2_in(n20805_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n20815_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n20816_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n20817_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n20818 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n20819 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n20820 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20815_o),
    .x1_in(n20816_o),
    .x2_in(n20817_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n20827_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n20828_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n20829_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n20830 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n20831 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n20832 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20827_o),
    .x1_in(n20828_o),
    .x2_in(n20829_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n20839_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n20840_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n20841_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n20842 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n20843 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n20844 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20839_o),
    .x1_in(n20840_o),
    .x2_in(n20841_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n20851_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n20852_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n20853_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n20854 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n20855 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n20856 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20851_o),
    .x1_in(n20852_o),
    .x2_in(n20853_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n20863_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n20864_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n20865_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n20866 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n20867 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n20868 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20863_o),
    .x1_in(n20864_o),
    .x2_in(n20865_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n20875_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n20876_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n20877_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n20878 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n20879 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n20880 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n20875_o),
    .x1_in(n20876_o),
    .x2_in(n20877_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n20887_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n20888_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n20889 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n20890 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n20891 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n20900 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n20901 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n20902_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n20903_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n20904 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n20905 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n20906 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n20907 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n20908 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n20909 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n20910 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n20911 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n20912 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n20913 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n20914 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n20915 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n20916 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n20902_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n20903_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n20949 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n20950 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n20951 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n20952 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n20953 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n20954 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n20955 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n20956 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n20957 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n20958 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n20959 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n20960 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n20961 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n20962 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n20963 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n20964 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n20965 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n20966 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n20967 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n20968 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n20969 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n20970 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n20971 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n20972 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n20973 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n20974 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n20975 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n20976 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n20977 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n20978 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_0_3 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n21039 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n21040 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n21041 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n21042 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n21043 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n21044 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n21045 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n21046 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n21047 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n21048 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n21049 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n21050 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n21051 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n21052 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n21053 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n21054 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n21055 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n21056 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n21057 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n21058 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n21059 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n21105_o = {alu_7_i_n20878, alu_6_i_n20866, alu_5_i_n20854, alu_4_i_n20842, alu_3_i_n20830, alu_2_i_n20818, alu_1_i_n20806, alu_0_i_n20794};
  assign n21106_o = {alu_7_i_n20880, alu_6_i_n20868, alu_5_i_n20856, alu_4_i_n20844, alu_3_i_n20832, alu_2_i_n20820, alu_1_i_n20808, alu_0_i_n20796};
  assign n21107_o = {alu_7_i_n20879, alu_6_i_n20867, alu_5_i_n20855, alu_4_i_n20843, alu_3_i_n20831, alu_2_i_n20819, alu_1_i_n20807, alu_0_i_n20795};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21108_o = dp_readena_vm ? n20670_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21109_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n21109_q <= n21108_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21110_o = dp_readena_vm ? n20671_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21111_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n21111_q <= n21110_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21112_q <= 1'b0;
    else
      n21112_q <= n20682_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21113_q <= 1'b0;
    else
      n21113_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21114_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21115_q <= 1'b0;
    else
      n21115_q <= n21114_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21116_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21117_q <= 2'b00;
    else
      n21117_q <= n21116_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21118_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21119_q <= 2'b00;
    else
      n21119_q <= n21118_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21120_o = dp_readena_vm ? n20675_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21121_q <= 3'b000;
    else
      n21121_q <= n21120_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21122_o = dp_readena_vm ? n20677_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21123_q <= 3'b000;
    else
      n21123_q <= n21122_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21124_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21125_q <= 1'b0;
    else
      n21125_q <= n21124_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n21126_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n20618_o)
    if (n20618_o)
      n21127_q <= 2'b00;
    else
      n21127_q <= n21126_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21128_q <= 3'b000;
    else
      n21128_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21129_q <= 3'b000;
    else
      n21129_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21130_q <= 2'b00;
    else
      n21130_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21133_q <= 3'b000;
    else
      n21133_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21134_q <= 3'b000;
    else
      n21134_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21135_q <= 1'b0;
    else
      n21135_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21136_q <= 2'b00;
    else
      n21136_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21137_q <= 2'b00;
    else
      n21137_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21138_q <= 1'b0;
    else
      n21138_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21139_q <= 2'b00;
    else
      n21139_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21140_q <= 22'b0000000000000000000000;
    else
      n21140_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21141_q <= 3'b000;
    else
      n21141_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21142_q <= 22'b0000000000000000000000;
    else
      n21142_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21143_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n21143_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21144_o = n20291_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21145_q <= 1'b0;
    else
      n21145_q <= n21144_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21146_o = n20291_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21147_q <= 1'b0;
    else
      n21147_q <= n21146_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21148_o = n20437_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21149_q <= 1'b0;
    else
      n21149_q <= n21148_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21152_q <= 22'b0000000000000000000000;
    else
      n21152_q <= n20289_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21153_q <= 22'b0000000000000000000000;
    else
      n21153_q <= n20435_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21154_o = n20437_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21155_q <= 6'b000000;
    else
      n21155_q <= n21154_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21156_o = n20437_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21157_q <= 1'b0;
    else
      n21157_q <= n21156_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21160_o = n20437_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21161_q <= 3'b000;
    else
      n21161_q <= n21160_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21162_o = n20437_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21163_q <= 2'b00;
    else
      n21163_q <= n21162_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21164_o = n20437_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21165_q <= 1'b0;
    else
      n21165_q <= n21164_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n21166_o = n20437_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21167_q <= 22'b0000000000000000000000;
    else
      n21167_q <= n21166_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21168_o = n20291_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21169_q <= 1'b0;
    else
      n21169_q <= n21168_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21170_o = n20291_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21171_q <= 3'b000;
    else
      n21171_q <= n21170_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21172_o = n20291_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21173_q <= 2'b00;
    else
      n21173_q <= n21172_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n21174_o = ~n20278_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n21175_o = n20291_o & n21174_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21176_o = n21175_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n21177_q <= n21176_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n21178_o = ~n20278_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n21179_o = n20291_o & n21178_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21180_o = n21179_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n21181_q <= n21180_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21182_o = n20291_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21183_q <= 1'b0;
    else
      n21183_q <= n21182_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21184_o = n20291_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21185_q <= 2'b00;
    else
      n21185_q <= n21184_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21186_o = n20291_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21187_q <= 2'b00;
    else
      n21187_q <= n21186_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21188_o = n20291_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21189_q <= 1'b0;
    else
      n21189_q <= n21188_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n21190_o = n20291_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21191_q <= 2'b00;
    else
      n21191_q <= n21190_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21192_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n21192_q <= n20449_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n21193_o = {n20492_o, n21192_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21194_q <= 3'b000;
    else
      n21194_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n20278_o)
    if (n20278_o)
      n21195_q <= 3'b000;
    else
      n21195_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n20424_o)
    if (n20424_o)
      n21196_q <= 3'b000;
    else
      n21196_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21198_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n21198_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21199_q <= 32'b00000000000000000000000000000000;
    else
      n21199_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21200_q <= 1'b0;
    else
      n21200_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21201_q <= 1'b0;
    else
      n21201_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21202_q <= 1'b0;
    else
      n21202_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21203_q <= 2'b00;
    else
      n21203_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21204_q <= 4'b0000;
    else
      n21204_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21205_q <= 1'b0;
    else
      n21205_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21206_q <= 4'b0000;
    else
      n21206_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21207_q <= 1'b0;
    else
      n21207_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21208_q <= 4'b0000;
    else
      n21208_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21209_q <= 1'b0;
    else
      n21209_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21210_q <= 1'b0;
    else
      n21210_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21211_q <= 2'b00;
    else
      n21211_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n20567_o)
    if (n20567_o)
      n21212_q <= 28'b0000000000000000000000000000;
    else
      n21212_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21213_q <= 1'b0;
    else
      n21213_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21214_q <= 1'b0;
    else
      n21214_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21216_q <= 1'b0;
    else
      n21216_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n20355_o)
    if (n20355_o)
      n21217_q <= 1'b0;
    else
      n21217_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21219_q <= 1'b0;
    else
      n21219_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21220_q <= 1'b0;
    else
      n21220_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21221_q <= 1'b0;
    else
      n21221_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21222_q <= 22'b0000000000000000000000;
    else
      n21222_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21223_q <= 1'b0;
    else
      n21223_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21224_q <= 22'b0000000000000000000000;
    else
      n21224_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21225_q <= 22'b0000000000000000000000;
    else
      n21225_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21226_q <= 1'b0;
    else
      n21226_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21227_q <= 22'b0000000000000000000000;
    else
      n21227_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21228_q <= 6'b000000;
    else
      n21228_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21229_q <= 1'b0;
    else
      n21229_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21230_q <= 1'b0;
    else
      n21230_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21231_q <= 1'b0;
    else
      n21231_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21232_q <= 3'b000;
    else
      n21232_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21233_q <= 2'b00;
    else
      n21233_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21234_q <= 1'b0;
    else
      n21234_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21235_q <= 1'b0;
    else
      n21235_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21236_q <= 3'b000;
    else
      n21236_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21237_q <= 2'b00;
    else
      n21237_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21238_q <= 1'b0;
    else
      n21238_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21239_q <= 2'b00;
    else
      n21239_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21240_q <= 2'b00;
    else
      n21240_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21241_q <= 1'b0;
    else
      n21241_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21242_q <= 2'b00;
    else
      n21242_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21243_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n21243_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n20082_o)
    if (n20082_o)
      n21244_q <= 1'b0;
    else
      n21244_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n21245_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n21246_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_0_2
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n18895_o;
  wire n18896_o;
  wire n18897_o;
  wire n18900_o;
  wire [4:0] n18988_o;
  wire n18989_o;
  wire [4:0] n18990_o;
  wire n18991_o;
  wire [2:0] n18994_o;
  wire [4:0] n18996_o;
  wire n18997_o;
  wire n18998_o;
  wire n18999_o;
  wire n19000_o;
  wire [4:0] n19001_o;
  wire [4:0] n19002_o;
  wire [4:0] n19003_o;
  wire n19004_o;
  wire n19005_o;
  wire n19006_o;
  wire [4:0] n19007_o;
  wire n19008_o;
  wire n19009_o;
  wire [4:0] n19010_o;
  wire n19011_o;
  wire n19012_o;
  wire n19013_o;
  wire n19014_o;
  wire n19017_o;
  wire n19023_o;
  wire n19025_o;
  wire [2:0] n19027_o;
  wire n19029_o;
  wire n19030_o;
  wire n19031_o;
  wire [2:0] n19033_o;
  wire [2:0] n19035_o;
  wire [2:0] n19037_o;
  wire n19038_o;
  wire n19039_o;
  wire [21:0] n19040_o;
  wire n19041_o;
  wire [2:0] n19042_o;
  wire [1:0] n19043_o;
  wire n19044_o;
  wire [21:0] n19045_o;
  wire n19046_o;
  wire [1:0] n19047_o;
  wire [1:0] n19048_o;
  wire n19049_o;
  wire [1:0] n19050_o;
  wire [2:0] n19051_o;
  wire [2:0] n19052_o;
  wire n19057_o;
  wire n19058_o;
  wire n19059_o;
  wire n19060_o;
  wire n19061_o;
  wire n19063_o;
  wire [2:0] n19065_o;
  wire n19067_o;
  wire n19068_o;
  wire n19069_o;
  wire [2:0] n19071_o;
  wire [2:0] n19075_o;
  wire [2:0] n19077_o;
  wire n19078_o;
  wire [21:0] n19080_o;
  wire [5:0] n19081_o;
  wire n19082_o;
  wire [2:0] n19083_o;
  wire [1:0] n19084_o;
  wire n19085_o;
  wire [21:0] n19086_o;
  wire [2:0] n19088_o;
  wire [2:0] n19091_o;
  wire n19096_o;
  wire n19099_o;
  wire n19100_o;
  wire [21:0] n19101_o;
  wire [21:0] n19103_o;
  wire [21:0] n19104_o;
  wire [21:0] n19106_o;
  wire [21:0] n19107_o;
  wire n19109_o;
  wire n19173_o;
  wire n19242_o;
  wire n19245_o;
  wire n19246_o;
  wire [21:0] n19247_o;
  wire [21:0] n19249_o;
  wire [21:0] n19250_o;
  wire [21:0] n19252_o;
  wire [21:0] n19253_o;
  wire n19255_o;
  wire [83:0] n19256_o;
  wire [83:0] n19257_o;
  wire [83:0] n19267_o;
  wire [11:0] n19309_o;
  wire [11:0] n19310_o;
  wire n19324_o;
  wire n19326_o;
  wire [11:0] n19327_o;
  wire [11:0] n19328_o;
  wire [11:0] n19329_o;
  wire [95:0] n19331_o;
  wire [95:0] n19332_o;
  wire [1:0] n19338_o;
  wire [2:0] n19339_o;
  wire n19340_o;
  wire n19342_o;
  wire n19343_o;
  wire n19345_o;
  wire n19346_o;
  wire n19349_o;
  wire n19351_o;
  wire n19352_o;
  wire n19355_o;
  wire n19356_o;
  wire [1:0] n19358_o;
  wire [1:0] n19360_o;
  wire n19362_o;
  wire [1:0] n19364_o;
  wire [1:0] n19370_o;
  wire [2:0] n19371_o;
  wire [4:0] n19372_o;
  wire n19375_o;
  wire [95:0] n19376_o;
  wire [95:0] n19378_o;
  wire n19380_o;
  wire n19385_o;
  wire n19436_o;
  wire n19439_o;
  wire [2:0] n19440_o;
  wire [11:0] n19441_o;
  wire n19443_o;
  wire [11:0] n19444_o;
  wire n19446_o;
  wire [11:0] n19447_o;
  wire n19449_o;
  wire [11:0] n19450_o;
  wire n19452_o;
  wire [11:0] n19453_o;
  wire n19455_o;
  wire [11:0] n19456_o;
  wire n19458_o;
  wire [11:0] n19459_o;
  wire n19461_o;
  wire [11:0] n19462_o;
  wire [6:0] n19463_o;
  wire [11:0] n19464_o;
  reg [11:0] n19465_o;
  wire [11:0] n19466_o;
  reg [11:0] n19467_o;
  wire [11:0] n19468_o;
  reg [11:0] n19469_o;
  wire [11:0] n19470_o;
  reg [11:0] n19471_o;
  wire [11:0] n19472_o;
  reg [11:0] n19473_o;
  wire [11:0] n19474_o;
  reg [11:0] n19475_o;
  wire [11:0] n19476_o;
  reg [11:0] n19477_o;
  wire [11:0] n19478_o;
  reg [11:0] n19479_o;
  wire n19481_o;
  wire n19484_o;
  wire [95:0] n19485_o;
  wire [95:0] n19486_o;
  wire [95:0] n19487_o;
  wire [95:0] n19488_o;
  wire [95:0] n19489_o;
  wire n19491_o;
  wire [2:0] n19493_o;
  wire [2:0] n19495_o;
  wire n19500_o;
  wire [12:0] xregister_file_i_n19549;
  wire [255:0] xregister_file_i_n19550;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n19555;
  wire [12:0] iregister_i_n19556;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n19563_o;
  wire n19565_o;
  wire n19566_o;
  wire n19568_o;
  wire n19569_o;
  wire n19572_o;
  wire n19574_o;
  wire n19575_o;
  wire n19578_o;
  wire n19579_o;
  wire [4:0] n19587_o;
  wire n19588_o;
  wire [4:0] n19589_o;
  wire [4:0] n19590_o;
  wire [4:0] n19592_o;
  wire n19593_o;
  wire n19594_o;
  wire n19595_o;
  wire n19597_o;
  wire n19598_o;
  wire n19600_o;
  wire n19601_o;
  wire n19602_o;
  wire n19603_o;
  wire n19606_o;
  wire [31:0] n19609_o;
  wire [11:0] n19610_o;
  wire [11:0] n19611_o;
  wire [31:0] alu_0_i_n19612;
  wire alu_0_i_n19613;
  wire [11:0] alu_0_i_n19614;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n19621_o;
  wire [11:0] n19622_o;
  wire [11:0] n19623_o;
  wire [31:0] alu_1_i_n19624;
  wire alu_1_i_n19625;
  wire [11:0] alu_1_i_n19626;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n19633_o;
  wire [11:0] n19634_o;
  wire [11:0] n19635_o;
  wire [31:0] alu_2_i_n19636;
  wire alu_2_i_n19637;
  wire [11:0] alu_2_i_n19638;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n19645_o;
  wire [11:0] n19646_o;
  wire [11:0] n19647_o;
  wire [31:0] alu_3_i_n19648;
  wire alu_3_i_n19649;
  wire [11:0] alu_3_i_n19650;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n19657_o;
  wire [11:0] n19658_o;
  wire [11:0] n19659_o;
  wire [31:0] alu_4_i_n19660;
  wire alu_4_i_n19661;
  wire [11:0] alu_4_i_n19662;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n19669_o;
  wire [11:0] n19670_o;
  wire [11:0] n19671_o;
  wire [31:0] alu_5_i_n19672;
  wire alu_5_i_n19673;
  wire [11:0] alu_5_i_n19674;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n19681_o;
  wire [11:0] n19682_o;
  wire [11:0] n19683_o;
  wire [31:0] alu_6_i_n19684;
  wire alu_6_i_n19685;
  wire [11:0] alu_6_i_n19686;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n19693_o;
  wire [11:0] n19694_o;
  wire [11:0] n19695_o;
  wire [31:0] alu_7_i_n19696;
  wire alu_7_i_n19697;
  wire [11:0] alu_7_i_n19698;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n19705_o;
  wire n19706_o;
  wire [12:0] ialu_i_n19707;
  wire ialu_i_n19708;
  wire ialu_i_n19709;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n19718;
  wire [95:0] register_bank_i_n19719;
  wire [16:0] n19720_o;
  wire [16:0] n19721_o;
  wire [95:0] register_bank_i_n19722;
  wire register_bank_i_n19723;
  wire register_bank_i_n19724;
  wire [2:0] register_bank_i_n19725;
  wire [2:0] register_bank_i_n19726;
  wire [1:0] register_bank_i_n19727;
  wire [2:0] register_bank_i_n19728;
  wire [2:0] register_bank_i_n19729;
  wire register_bank_i_n19730;
  wire [1:0] register_bank_i_n19731;
  wire [1:0] register_bank_i_n19732;
  wire register_bank_i_n19733;
  wire [1:0] register_bank_i_n19734;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n19767;
  wire instr_decoder2_i_n19768;
  wire [3:0] instr_decoder2_i_n19769;
  wire instr_decoder2_i_n19770;
  wire instr_decoder2_i_n19771;
  wire instr_decoder2_i_n19772;
  wire instr_decoder2_i_n19773;
  wire [11:0] instr_decoder2_i_n19774;
  wire [11:0] instr_decoder2_i_n19775;
  wire [11:0] instr_decoder2_i_n19776;
  wire instr_decoder2_i_n19777;
  wire instr_decoder2_i_n19778;
  wire instr_decoder2_i_n19779;
  wire [7:0] instr_decoder2_i_n19780;
  wire instr_decoder2_i_n19781;
  wire [11:0] instr_decoder2_i_n19782;
  wire instr_decoder2_i_n19783;
  wire instr_decoder2_i_n19784;
  wire [3:0] instr_decoder2_i_n19785;
  wire [3:0] instr_decoder2_i_n19786;
  wire instr_decoder2_i_n19787;
  wire instr_decoder2_i_n19788;
  wire [2:0] instr_decoder2_i_n19789;
  wire [12:0] instr_decoder2_i_n19790;
  wire instr_decoder2_i_n19791;
  wire [4:0] instr_decoder2_i_n19792;
  wire [12:0] instr_decoder2_i_n19793;
  wire [12:0] instr_decoder2_i_n19794;
  wire [7:0] instr_decoder2_i_n19795;
  wire [7:0] instr_decoder2_i_n19796;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n19857;
  wire instr_dispatch2_i1_n19858;
  wire [11:0] instr_dispatch2_i1_n19859;
  wire [11:0] instr_dispatch2_i1_n19860;
  wire instr_dispatch2_i1_n19861;
  wire instr_dispatch2_i1_n19862;
  wire instr_dispatch2_i1_n19863;
  wire instr_dispatch2_i1_n19864;
  wire instr_dispatch2_i1_n19865;
  wire instr_dispatch2_i1_n19866;
  wire instr_dispatch2_i1_n19867;
  wire instr_dispatch2_i1_n19868;
  wire [11:0] instr_dispatch2_i1_n19869;
  wire [7:0] instr_dispatch2_i1_n19870;
  wire [95:0] instr_dispatch2_i1_n19871;
  wire [7:0] instr_dispatch2_i1_n19872;
  wire [95:0] instr_dispatch2_i1_n19873;
  wire [95:0] instr_dispatch2_i1_n19874;
  wire [11:0] instr_dispatch2_i1_n19875;
  wire [4:0] instr_dispatch2_i1_n19876;
  wire [3:0] instr_dispatch2_i1_n19877;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n19923_o;
  wire [95:0] n19924_o;
  wire [7:0] n19925_o;
  wire [95:0] n19926_o;
  reg [95:0] n19927_q;
  wire [95:0] n19928_o;
  reg [95:0] n19929_q;
  reg n19930_q;
  reg n19931_q;
  wire n19932_o;
  reg n19933_q;
  wire [1:0] n19934_o;
  reg [1:0] n19935_q;
  wire [1:0] n19936_o;
  reg [1:0] n19937_q;
  wire [2:0] n19938_o;
  reg [2:0] n19939_q;
  wire [2:0] n19940_o;
  reg [2:0] n19941_q;
  wire n19942_o;
  reg n19943_q;
  wire [1:0] n19944_o;
  reg [1:0] n19945_q;
  reg [2:0] n19946_q;
  reg [2:0] n19947_q;
  reg [1:0] n19948_q;
  reg [2:0] n19951_q;
  reg [2:0] n19952_q;
  reg n19953_q;
  reg [1:0] n19954_q;
  reg [1:0] n19955_q;
  reg n19956_q;
  reg [1:0] n19957_q;
  reg [21:0] n19958_q;
  reg [2:0] n19959_q;
  reg [21:0] n19960_q;
  reg [95:0] n19961_q;
  wire n19962_o;
  reg n19963_q;
  wire n19964_o;
  reg n19965_q;
  wire n19966_o;
  reg n19967_q;
  reg [21:0] n19970_q;
  reg [21:0] n19971_q;
  wire [5:0] n19972_o;
  reg [5:0] n19973_q;
  wire n19974_o;
  reg n19975_q;
  wire [2:0] n19978_o;
  reg [2:0] n19979_q;
  wire [1:0] n19980_o;
  reg [1:0] n19981_q;
  wire n19982_o;
  reg n19983_q;
  wire [21:0] n19984_o;
  reg [21:0] n19985_q;
  wire n19986_o;
  reg n19987_q;
  wire [2:0] n19988_o;
  reg [2:0] n19989_q;
  wire [1:0] n19990_o;
  reg [1:0] n19991_q;
  wire n19992_o;
  wire n19993_o;
  wire n19994_o;
  reg n19995_q;
  wire n19996_o;
  wire n19997_o;
  wire [21:0] n19998_o;
  reg [21:0] n19999_q;
  wire n20000_o;
  reg n20001_q;
  wire [1:0] n20002_o;
  reg [1:0] n20003_q;
  wire [1:0] n20004_o;
  reg [1:0] n20005_q;
  wire n20006_o;
  reg n20007_q;
  wire [1:0] n20008_o;
  reg [1:0] n20009_q;
  reg [83:0] n20010_q;
  wire [95:0] n20011_o;
  reg [2:0] n20012_q;
  reg [2:0] n20013_q;
  reg [2:0] n20014_q;
  reg [79:0] n20016_q;
  reg [31:0] n20017_q;
  reg n20018_q;
  reg n20019_q;
  reg n20020_q;
  reg [1:0] n20021_q;
  reg [3:0] n20022_q;
  reg n20023_q;
  reg [3:0] n20024_q;
  reg n20025_q;
  reg [3:0] n20026_q;
  reg n20027_q;
  reg n20028_q;
  reg [1:0] n20029_q;
  reg [27:0] n20030_q;
  reg n20031_q;
  reg n20032_q;
  reg n20034_q;
  reg n20035_q;
  reg n20037_q;
  reg n20038_q;
  reg n20039_q;
  reg [21:0] n20040_q;
  reg n20041_q;
  reg [21:0] n20042_q;
  reg [21:0] n20043_q;
  reg n20044_q;
  reg [21:0] n20045_q;
  reg [5:0] n20046_q;
  reg n20047_q;
  reg n20048_q;
  reg n20049_q;
  reg [2:0] n20050_q;
  reg [1:0] n20051_q;
  reg n20052_q;
  reg n20053_q;
  reg [2:0] n20054_q;
  reg [1:0] n20055_q;
  reg n20056_q;
  reg [1:0] n20057_q;
  reg [1:0] n20058_q;
  reg n20059_q;
  reg [1:0] n20060_q;
  reg [95:0] n20061_q;
  reg n20062_q;
  wire [2:0] n20063_o;
  wire [2:0] n20064_o;
  assign i_y_neg_out = n19705_o;
  assign i_y_zero_out = n19706_o;
  assign dp_readdata_out = n19378_o;
  assign dp_readdata_vm_out = n19380_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n20063_o;
  assign dp_read_vaddr_out = n20064_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n19358_o;
  assign dp_read_data_type_out = n19360_o;
  assign dp_read_stream_out = n19362_o;
  assign dp_read_stream_id_out = n19364_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n19718; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n19719; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n19857; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n19858; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n19866; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n19863; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n19864; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n19865; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n19871; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n19872; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n19774; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n19775; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n19776; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n19556; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n19791; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n19767; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n19873; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n19874; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n19875; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n19923_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n19924_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n19925_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n19876; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n19877; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n19769; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n19606_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n19579_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n19372_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n19859; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n19860; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n19869; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n19870; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n19370_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n19371_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n19768; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n19773; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n19770; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n19771; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n19772; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n19781; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n19782; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n19777; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n19778; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n19779; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n19780; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n19861; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n19862; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n19868; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n19783; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n19784; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n19785; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n19555; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n19786; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n19787; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n19788; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n19789; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n19790; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n19927_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n19929_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n19930_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n19931_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n19933_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n19935_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n19937_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n19939_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n19941_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n19943_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n19945_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n19792; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n19793; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n19794; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n19707; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n19708; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n19709; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n19867; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n19795; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n19796; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n19549; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n19550; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n19038_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n19039_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n19078_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n19040_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n19080_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n19081_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n19082_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n19083_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n19084_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n19085_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n19086_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n19041_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n19042_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n19043_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n19044_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n19045_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n19046_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n19047_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n19048_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n19049_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n19050_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n19332_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n19051_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n19052_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n19088_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n19091_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n19946_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n19947_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n19948_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n19951_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n19952_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n19953_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n19954_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n19955_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n19956_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n19957_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n19958_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n19959_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n19960_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n19961_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n19963_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n19965_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n19967_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n19970_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n19971_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n19973_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n19975_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n19979_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n19981_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n19983_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n19985_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n19987_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n19989_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n19991_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n19995_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n19999_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n20001_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n20003_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n20005_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n20007_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n20009_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n20011_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n20012_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n20013_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n20014_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n19356_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n19017_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n19724; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n19725; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n19726; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n19727; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n19728; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n19729; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n19722; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n19723; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n19730; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n19731; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n19732; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n19733; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n19734; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n18895_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n18896_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n18897_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n20016_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n20017_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n20018_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n20019_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n20020_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n20021_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n20022_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n20023_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n20024_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n20025_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n20026_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n20027_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n20028_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n20029_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n20030_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n20031_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n20032_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n20034_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n20035_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n20037_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n20038_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n20039_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n20040_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n20041_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n20042_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n20043_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n20044_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n20045_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n20046_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n20047_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n20048_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n20049_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n20050_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n20051_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n20052_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n20053_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n20054_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n20055_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n20056_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n20057_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n20058_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n20059_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n20060_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n20061_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n20062_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n18895_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n18896_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n18897_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n18900_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n18988_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n18989_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n18990_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n18991_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n18994_o = n18991_o ? 3'b000 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n18996_o = n18990_o + n18988_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n18997_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n18998_o = n18997_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n18999_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n19000_o = n18999_o & n18998_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n19001_o = n18988_o & n18990_o;
  /* ../../HW/src/pcore/pcore.vhd:215:8  */
  assign n19002_o = {n18994_o, 2'b10};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n19003_o = n18988_o & n19002_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n19004_o = n19001_o == n19003_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n19005_o = n19004_o & n18989_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n19006_o = ~n18989_o;
  /* ../../HW/src/pcore/pcore.vhd:106:8  */
  assign n19007_o = {n18994_o, 2'b10};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n19008_o = $unsigned(n19007_o) >= $unsigned(n18990_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n19009_o = n19008_o & n19006_o;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n19010_o = {n18994_o, 2'b10};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n19011_o = $unsigned(n19010_o) <= $unsigned(n18996_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n19012_o = n19011_o & n19009_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n19013_o = n19005_o | n19012_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n19014_o = n19013_o & n19000_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n19017_o = n19014_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n19023_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n19025_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n19027_o = n19025_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n19029_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n19030_o = n19029_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n19031_o = dp_read_gen_valid_in_r & n19030_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n19033_o = n19031_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n19035_o = n19031_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n19037_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19038_o = n19023_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19039_o = n19023_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19040_o = n19023_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19041_o = n19023_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19042_o = n19023_o ? n19027_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19043_o = n19023_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19044_o = n19023_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19045_o = n19023_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19046_o = n19023_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19047_o = n19023_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19048_o = n19023_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19049_o = n19023_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19050_o = n19023_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19051_o = n19023_o ? n19033_o : n19037_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n19052_o = n19023_o ? n19035_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n19057_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n19058_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n19059_o = dp_write_in_r & n19058_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n19060_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n19061_o = n19059_o & n19060_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n19063_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n19065_o = n19063_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n19067_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n19068_o = n19067_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n19069_o = dp_write_gen_valid_in_r & n19068_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n19071_o = n19069_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n19075_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n19077_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19078_o = n19057_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19080_o = n19057_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19081_o = n19057_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19082_o = n19057_o ? n19061_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19083_o = n19057_o ? n19065_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19084_o = n19057_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19085_o = n19057_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19086_o = n19057_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19088_o = n19057_o ? n19071_o : n19075_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n19091_o = n19057_o ? 3'b000 : n19077_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n19096_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n19099_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n19100_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n19101_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n19103_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n19104_o = n19100_o ? n19101_o : n19103_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n19106_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n19107_o = n19099_o ? n19104_o : n19106_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n19109_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n19173_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n19242_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n19245_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n19246_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n19247_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n19249_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n19250_o = n19246_o ? n19247_o : n19249_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n19252_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n19253_o = n19245_o ? n19250_o : n19252_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n19255_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n19256_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n19257_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n19267_o = n19255_o ? n19256_o : n19257_o;
  assign n19309_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n19310_o = n19242_o ? 12'b000000000000 : n19309_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n19324_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n19326_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n19327_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n19328_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n19329_o = n19326_o ? n19327_o : n19328_o;
  assign n19331_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n19329_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n19332_o = n19324_o ? n19331_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n19338_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n19339_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n19340_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n19342_o = n19338_o == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n19343_o = n19342_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n19345_o = n19339_o == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n19346_o = n19345_o & n19343_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n19349_o = n19346_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n19351_o = n19338_o == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n19352_o = n19351_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n19355_o = n19352_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n19356_o = n19340_o ? n19349_o : n19355_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n19358_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n19360_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n19362_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n19364_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n19370_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n19371_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n19372_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n19375_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n19376_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n19378_o = n19375_o ? 96'bZ : n19376_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n19380_o = n19375_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n19385_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n19436_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n19439_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n19440_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n19441_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n19443_o = n19440_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n19444_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n19446_o = n19440_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n19447_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n19449_o = n19440_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n19450_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n19452_o = n19440_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n19453_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n19455_o = n19440_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n19456_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n19458_o = n19440_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n19459_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n19461_o = n19440_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n19462_o = dp_readdata_vm[11:0];
  assign n19463_o = {n19461_o, n19458_o, n19455_o, n19452_o, n19449_o, n19446_o, n19443_o};
  assign n19464_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19465_o = n19464_o;
      7'b0100000: n19465_o = n19464_o;
      7'b0010000: n19465_o = n19464_o;
      7'b0001000: n19465_o = n19464_o;
      7'b0000100: n19465_o = n19464_o;
      7'b0000010: n19465_o = n19464_o;
      7'b0000001: n19465_o = n19464_o;
      default: n19465_o = n19462_o;
    endcase
  assign n19466_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19467_o = n19459_o;
      7'b0100000: n19467_o = n19466_o;
      7'b0010000: n19467_o = n19466_o;
      7'b0001000: n19467_o = n19466_o;
      7'b0000100: n19467_o = n19466_o;
      7'b0000010: n19467_o = n19466_o;
      7'b0000001: n19467_o = n19466_o;
      default: n19467_o = n19466_o;
    endcase
  assign n19468_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19469_o = n19468_o;
      7'b0100000: n19469_o = n19456_o;
      7'b0010000: n19469_o = n19468_o;
      7'b0001000: n19469_o = n19468_o;
      7'b0000100: n19469_o = n19468_o;
      7'b0000010: n19469_o = n19468_o;
      7'b0000001: n19469_o = n19468_o;
      default: n19469_o = n19468_o;
    endcase
  assign n19470_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19471_o = n19470_o;
      7'b0100000: n19471_o = n19470_o;
      7'b0010000: n19471_o = n19453_o;
      7'b0001000: n19471_o = n19470_o;
      7'b0000100: n19471_o = n19470_o;
      7'b0000010: n19471_o = n19470_o;
      7'b0000001: n19471_o = n19470_o;
      default: n19471_o = n19470_o;
    endcase
  assign n19472_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19473_o = n19472_o;
      7'b0100000: n19473_o = n19472_o;
      7'b0010000: n19473_o = n19472_o;
      7'b0001000: n19473_o = n19450_o;
      7'b0000100: n19473_o = n19472_o;
      7'b0000010: n19473_o = n19472_o;
      7'b0000001: n19473_o = n19472_o;
      default: n19473_o = n19472_o;
    endcase
  assign n19474_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19475_o = n19474_o;
      7'b0100000: n19475_o = n19474_o;
      7'b0010000: n19475_o = n19474_o;
      7'b0001000: n19475_o = n19474_o;
      7'b0000100: n19475_o = n19447_o;
      7'b0000010: n19475_o = n19474_o;
      7'b0000001: n19475_o = n19474_o;
      default: n19475_o = n19474_o;
    endcase
  assign n19476_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19477_o = n19476_o;
      7'b0100000: n19477_o = n19476_o;
      7'b0010000: n19477_o = n19476_o;
      7'b0001000: n19477_o = n19476_o;
      7'b0000100: n19477_o = n19476_o;
      7'b0000010: n19477_o = n19444_o;
      7'b0000001: n19477_o = n19476_o;
      default: n19477_o = n19476_o;
    endcase
  assign n19478_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n19463_o)
      7'b1000000: n19479_o = n19478_o;
      7'b0100000: n19479_o = n19478_o;
      7'b0010000: n19479_o = n19478_o;
      7'b0001000: n19479_o = n19478_o;
      7'b0000100: n19479_o = n19478_o;
      7'b0000010: n19479_o = n19478_o;
      7'b0000001: n19479_o = n19441_o;
      default: n19479_o = n19478_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n19481_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n19484_o = n19481_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n19485_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n19486_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n19487_o = {n19479_o, n19477_o, n19475_o, n19473_o, n19471_o, n19469_o, n19467_o, n19465_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n19488_o = n19439_o ? n19487_o : n19485_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n19489_o = n19439_o ? dp_readdata2_r : n19486_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n19491_o = n19439_o ? n19484_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n19493_o = n19439_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n19495_o = n19439_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n19500_o = dp_readena_vm ? n19491_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n19549 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n19550 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n19555 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n19556 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n19563_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n19565_o = dp_rd_pid == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n19566_o = n19565_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n19568_o = dp_rd_cid == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n19569_o = n19568_o & n19566_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n19572_o = n19569_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n19574_o = dp_rd_pid == 2'b10;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n19575_o = n19574_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n19578_o = n19575_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n19579_o = n19563_o ? n19572_o : n19578_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n19587_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n19588_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n19589_o = dp_mcast_addr + n19587_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n19590_o = n19587_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n19592_o = n19587_o & 5'b00010;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n19593_o = n19590_o == n19592_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n19594_o = n19593_o & n19588_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n19595_o = ~n19588_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n19597_o = $unsigned(5'b00010) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n19598_o = n19597_o & n19595_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n19600_o = $unsigned(5'b00010) <= $unsigned(n19589_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n19601_o = n19600_o & n19598_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n19602_o = n19594_o | n19601_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n19603_o = n19602_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n19606_o = n19603_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n19609_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n19610_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n19611_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n19612 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n19613 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n19614 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19609_o),
    .x1_in(n19610_o),
    .x2_in(n19611_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n19621_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n19622_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n19623_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n19624 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n19625 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n19626 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19621_o),
    .x1_in(n19622_o),
    .x2_in(n19623_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n19633_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n19634_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n19635_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n19636 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n19637 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n19638 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19633_o),
    .x1_in(n19634_o),
    .x2_in(n19635_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n19645_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n19646_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n19647_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n19648 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n19649 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n19650 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19645_o),
    .x1_in(n19646_o),
    .x2_in(n19647_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n19657_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n19658_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n19659_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n19660 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n19661 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n19662 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19657_o),
    .x1_in(n19658_o),
    .x2_in(n19659_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n19669_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n19670_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n19671_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n19672 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n19673 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n19674 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19669_o),
    .x1_in(n19670_o),
    .x2_in(n19671_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n19681_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n19682_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n19683_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n19684 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n19685 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n19686 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19681_o),
    .x1_in(n19682_o),
    .x2_in(n19683_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n19693_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n19694_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n19695_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n19696 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n19697 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n19698 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n19693_o),
    .x1_in(n19694_o),
    .x2_in(n19695_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n19705_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n19706_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n19707 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n19708 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n19709 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n19718 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n19719 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n19720_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n19721_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n19722 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n19723 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n19724 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n19725 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n19726 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n19727 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n19728 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n19729 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n19730 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n19731 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n19732 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n19733 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n19734 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n19720_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n19721_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n19767 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n19768 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n19769 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n19770 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n19771 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n19772 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n19773 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n19774 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n19775 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n19776 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n19777 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n19778 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n19779 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n19780 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n19781 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n19782 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n19783 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n19784 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n19785 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n19786 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n19787 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n19788 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n19789 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n19790 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n19791 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n19792 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n19793 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n19794 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n19795 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n19796 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_0_2 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n19857 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n19858 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n19859 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n19860 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n19861 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n19862 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n19863 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n19864 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n19865 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n19866 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n19867 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n19868 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n19869 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n19870 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n19871 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n19872 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n19873 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n19874 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n19875 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n19876 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n19877 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n19923_o = {alu_7_i_n19696, alu_6_i_n19684, alu_5_i_n19672, alu_4_i_n19660, alu_3_i_n19648, alu_2_i_n19636, alu_1_i_n19624, alu_0_i_n19612};
  assign n19924_o = {alu_7_i_n19698, alu_6_i_n19686, alu_5_i_n19674, alu_4_i_n19662, alu_3_i_n19650, alu_2_i_n19638, alu_1_i_n19626, alu_0_i_n19614};
  assign n19925_o = {alu_7_i_n19697, alu_6_i_n19685, alu_5_i_n19673, alu_4_i_n19661, alu_3_i_n19649, alu_2_i_n19637, alu_1_i_n19625, alu_0_i_n19613};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19926_o = dp_readena_vm ? n19488_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19927_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n19927_q <= n19926_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19928_o = dp_readena_vm ? n19489_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19929_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n19929_q <= n19928_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19930_q <= 1'b0;
    else
      n19930_q <= n19500_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19931_q <= 1'b0;
    else
      n19931_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19932_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19933_q <= 1'b0;
    else
      n19933_q <= n19932_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19934_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19935_q <= 2'b00;
    else
      n19935_q <= n19934_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19936_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19937_q <= 2'b00;
    else
      n19937_q <= n19936_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19938_o = dp_readena_vm ? n19493_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19939_q <= 3'b000;
    else
      n19939_q <= n19938_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19940_o = dp_readena_vm ? n19495_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19941_q <= 3'b000;
    else
      n19941_q <= n19940_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19942_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19943_q <= 1'b0;
    else
      n19943_q <= n19942_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n19944_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n19436_o)
    if (n19436_o)
      n19945_q <= 2'b00;
    else
      n19945_q <= n19944_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19946_q <= 3'b000;
    else
      n19946_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19947_q <= 3'b000;
    else
      n19947_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19948_q <= 2'b00;
    else
      n19948_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19951_q <= 3'b000;
    else
      n19951_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19952_q <= 3'b000;
    else
      n19952_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19953_q <= 1'b0;
    else
      n19953_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19954_q <= 2'b00;
    else
      n19954_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19955_q <= 2'b00;
    else
      n19955_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19956_q <= 1'b0;
    else
      n19956_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19957_q <= 2'b00;
    else
      n19957_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19958_q <= 22'b0000000000000000000000;
    else
      n19958_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19959_q <= 3'b000;
    else
      n19959_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19960_q <= 22'b0000000000000000000000;
    else
      n19960_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n19961_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n19961_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19962_o = n19109_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n19963_q <= 1'b0;
    else
      n19963_q <= n19962_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19964_o = n19109_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n19965_q <= 1'b0;
    else
      n19965_q <= n19964_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19966_o = n19255_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19967_q <= 1'b0;
    else
      n19967_q <= n19966_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n19970_q <= 22'b0000000000000000000000;
    else
      n19970_q <= n19107_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19971_q <= 22'b0000000000000000000000;
    else
      n19971_q <= n19253_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19972_o = n19255_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19973_q <= 6'b000000;
    else
      n19973_q <= n19972_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19974_o = n19255_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19975_q <= 1'b0;
    else
      n19975_q <= n19974_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19978_o = n19255_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19979_q <= 3'b000;
    else
      n19979_q <= n19978_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19980_o = n19255_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19981_q <= 2'b00;
    else
      n19981_q <= n19980_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19982_o = n19255_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19983_q <= 1'b0;
    else
      n19983_q <= n19982_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n19984_o = n19255_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n19985_q <= 22'b0000000000000000000000;
    else
      n19985_q <= n19984_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19986_o = n19109_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n19987_q <= 1'b0;
    else
      n19987_q <= n19986_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19988_o = n19109_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n19989_q <= 3'b000;
    else
      n19989_q <= n19988_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19990_o = n19109_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n19991_q <= 2'b00;
    else
      n19991_q <= n19990_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n19992_o = ~n19096_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n19993_o = n19109_o & n19992_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19994_o = n19993_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n19995_q <= n19994_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n19996_o = ~n19096_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n19997_o = n19109_o & n19996_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n19998_o = n19997_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n19999_q <= n19998_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n20000_o = n19109_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20001_q <= 1'b0;
    else
      n20001_q <= n20000_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n20002_o = n19109_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20003_q <= 2'b00;
    else
      n20003_q <= n20002_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n20004_o = n19109_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20005_q <= 2'b00;
    else
      n20005_q <= n20004_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n20006_o = n19109_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20007_q <= 1'b0;
    else
      n20007_q <= n20006_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n20008_o = n19109_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20009_q <= 2'b00;
    else
      n20009_q <= n20008_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n20010_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n20010_q <= n19267_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n20011_o = {n19310_o, n20010_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20012_q <= 3'b000;
    else
      n20012_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n19096_o)
    if (n19096_o)
      n20013_q <= 3'b000;
    else
      n20013_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n19242_o)
    if (n19242_o)
      n20014_q <= 3'b000;
    else
      n20014_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20016_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n20016_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20017_q <= 32'b00000000000000000000000000000000;
    else
      n20017_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20018_q <= 1'b0;
    else
      n20018_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20019_q <= 1'b0;
    else
      n20019_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20020_q <= 1'b0;
    else
      n20020_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20021_q <= 2'b00;
    else
      n20021_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20022_q <= 4'b0000;
    else
      n20022_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20023_q <= 1'b0;
    else
      n20023_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20024_q <= 4'b0000;
    else
      n20024_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20025_q <= 1'b0;
    else
      n20025_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20026_q <= 4'b0000;
    else
      n20026_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20027_q <= 1'b0;
    else
      n20027_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20028_q <= 1'b0;
    else
      n20028_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20029_q <= 2'b00;
    else
      n20029_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n19385_o)
    if (n19385_o)
      n20030_q <= 28'b0000000000000000000000000000;
    else
      n20030_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n20031_q <= 1'b0;
    else
      n20031_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n20032_q <= 1'b0;
    else
      n20032_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n20034_q <= 1'b0;
    else
      n20034_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n19173_o)
    if (n19173_o)
      n20035_q <= 1'b0;
    else
      n20035_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20037_q <= 1'b0;
    else
      n20037_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20038_q <= 1'b0;
    else
      n20038_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20039_q <= 1'b0;
    else
      n20039_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20040_q <= 22'b0000000000000000000000;
    else
      n20040_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20041_q <= 1'b0;
    else
      n20041_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20042_q <= 22'b0000000000000000000000;
    else
      n20042_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20043_q <= 22'b0000000000000000000000;
    else
      n20043_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20044_q <= 1'b0;
    else
      n20044_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20045_q <= 22'b0000000000000000000000;
    else
      n20045_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20046_q <= 6'b000000;
    else
      n20046_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20047_q <= 1'b0;
    else
      n20047_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20048_q <= 1'b0;
    else
      n20048_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20049_q <= 1'b0;
    else
      n20049_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20050_q <= 3'b000;
    else
      n20050_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20051_q <= 2'b00;
    else
      n20051_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20052_q <= 1'b0;
    else
      n20052_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20053_q <= 1'b0;
    else
      n20053_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20054_q <= 3'b000;
    else
      n20054_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20055_q <= 2'b00;
    else
      n20055_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20056_q <= 1'b0;
    else
      n20056_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20057_q <= 2'b00;
    else
      n20057_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20058_q <= 2'b00;
    else
      n20058_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20059_q <= 1'b0;
    else
      n20059_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20060_q <= 2'b00;
    else
      n20060_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20061_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n20061_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n18900_o)
    if (n18900_o)
      n20062_q <= 1'b0;
    else
      n20062_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n20063_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n20064_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_0_1
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n17713_o;
  wire n17714_o;
  wire n17715_o;
  wire n17718_o;
  wire [4:0] n17806_o;
  wire n17807_o;
  wire [4:0] n17808_o;
  wire n17809_o;
  wire [2:0] n17812_o;
  wire [4:0] n17814_o;
  wire n17815_o;
  wire n17816_o;
  wire n17817_o;
  wire n17818_o;
  wire [4:0] n17819_o;
  wire [4:0] n17820_o;
  wire [4:0] n17821_o;
  wire n17822_o;
  wire n17823_o;
  wire n17824_o;
  wire [4:0] n17825_o;
  wire n17826_o;
  wire n17827_o;
  wire [4:0] n17828_o;
  wire n17829_o;
  wire n17830_o;
  wire n17831_o;
  wire n17832_o;
  wire n17835_o;
  wire n17841_o;
  wire n17843_o;
  wire [2:0] n17845_o;
  wire n17847_o;
  wire n17848_o;
  wire n17849_o;
  wire [2:0] n17851_o;
  wire [2:0] n17853_o;
  wire [2:0] n17855_o;
  wire n17856_o;
  wire n17857_o;
  wire [21:0] n17858_o;
  wire n17859_o;
  wire [2:0] n17860_o;
  wire [1:0] n17861_o;
  wire n17862_o;
  wire [21:0] n17863_o;
  wire n17864_o;
  wire [1:0] n17865_o;
  wire [1:0] n17866_o;
  wire n17867_o;
  wire [1:0] n17868_o;
  wire [2:0] n17869_o;
  wire [2:0] n17870_o;
  wire n17875_o;
  wire n17876_o;
  wire n17877_o;
  wire n17878_o;
  wire n17879_o;
  wire n17881_o;
  wire [2:0] n17883_o;
  wire n17885_o;
  wire n17886_o;
  wire n17887_o;
  wire [2:0] n17889_o;
  wire [2:0] n17893_o;
  wire [2:0] n17895_o;
  wire n17896_o;
  wire [21:0] n17898_o;
  wire [5:0] n17899_o;
  wire n17900_o;
  wire [2:0] n17901_o;
  wire [1:0] n17902_o;
  wire n17903_o;
  wire [21:0] n17904_o;
  wire [2:0] n17906_o;
  wire [2:0] n17909_o;
  wire n17914_o;
  wire n17917_o;
  wire n17918_o;
  wire [21:0] n17919_o;
  wire [21:0] n17921_o;
  wire [21:0] n17922_o;
  wire [21:0] n17924_o;
  wire [21:0] n17925_o;
  wire n17927_o;
  wire n17991_o;
  wire n18060_o;
  wire n18063_o;
  wire n18064_o;
  wire [21:0] n18065_o;
  wire [21:0] n18067_o;
  wire [21:0] n18068_o;
  wire [21:0] n18070_o;
  wire [21:0] n18071_o;
  wire n18073_o;
  wire [83:0] n18074_o;
  wire [83:0] n18075_o;
  wire [83:0] n18085_o;
  wire [11:0] n18127_o;
  wire [11:0] n18128_o;
  wire n18142_o;
  wire n18144_o;
  wire [11:0] n18145_o;
  wire [11:0] n18146_o;
  wire [11:0] n18147_o;
  wire [95:0] n18149_o;
  wire [95:0] n18150_o;
  wire [1:0] n18156_o;
  wire [2:0] n18157_o;
  wire n18158_o;
  wire n18160_o;
  wire n18161_o;
  wire n18163_o;
  wire n18164_o;
  wire n18167_o;
  wire n18169_o;
  wire n18170_o;
  wire n18173_o;
  wire n18174_o;
  wire [1:0] n18176_o;
  wire [1:0] n18178_o;
  wire n18180_o;
  wire [1:0] n18182_o;
  wire [1:0] n18188_o;
  wire [2:0] n18189_o;
  wire [4:0] n18190_o;
  wire n18193_o;
  wire [95:0] n18194_o;
  wire [95:0] n18196_o;
  wire n18198_o;
  wire n18203_o;
  wire n18254_o;
  wire n18257_o;
  wire [2:0] n18258_o;
  wire [11:0] n18259_o;
  wire n18261_o;
  wire [11:0] n18262_o;
  wire n18264_o;
  wire [11:0] n18265_o;
  wire n18267_o;
  wire [11:0] n18268_o;
  wire n18270_o;
  wire [11:0] n18271_o;
  wire n18273_o;
  wire [11:0] n18274_o;
  wire n18276_o;
  wire [11:0] n18277_o;
  wire n18279_o;
  wire [11:0] n18280_o;
  wire [6:0] n18281_o;
  wire [11:0] n18282_o;
  reg [11:0] n18283_o;
  wire [11:0] n18284_o;
  reg [11:0] n18285_o;
  wire [11:0] n18286_o;
  reg [11:0] n18287_o;
  wire [11:0] n18288_o;
  reg [11:0] n18289_o;
  wire [11:0] n18290_o;
  reg [11:0] n18291_o;
  wire [11:0] n18292_o;
  reg [11:0] n18293_o;
  wire [11:0] n18294_o;
  reg [11:0] n18295_o;
  wire [11:0] n18296_o;
  reg [11:0] n18297_o;
  wire n18299_o;
  wire n18302_o;
  wire [95:0] n18303_o;
  wire [95:0] n18304_o;
  wire [95:0] n18305_o;
  wire [95:0] n18306_o;
  wire [95:0] n18307_o;
  wire n18309_o;
  wire [2:0] n18311_o;
  wire [2:0] n18313_o;
  wire n18318_o;
  wire [12:0] xregister_file_i_n18367;
  wire [255:0] xregister_file_i_n18368;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n18373;
  wire [12:0] iregister_i_n18374;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n18381_o;
  wire n18383_o;
  wire n18384_o;
  wire n18386_o;
  wire n18387_o;
  wire n18390_o;
  wire n18392_o;
  wire n18393_o;
  wire n18396_o;
  wire n18397_o;
  wire [4:0] n18405_o;
  wire n18406_o;
  wire [4:0] n18407_o;
  wire [4:0] n18408_o;
  wire [4:0] n18410_o;
  wire n18411_o;
  wire n18412_o;
  wire n18413_o;
  wire n18415_o;
  wire n18416_o;
  wire n18418_o;
  wire n18419_o;
  wire n18420_o;
  wire n18421_o;
  wire n18424_o;
  wire [31:0] n18427_o;
  wire [11:0] n18428_o;
  wire [11:0] n18429_o;
  wire [31:0] alu_0_i_n18430;
  wire alu_0_i_n18431;
  wire [11:0] alu_0_i_n18432;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n18439_o;
  wire [11:0] n18440_o;
  wire [11:0] n18441_o;
  wire [31:0] alu_1_i_n18442;
  wire alu_1_i_n18443;
  wire [11:0] alu_1_i_n18444;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n18451_o;
  wire [11:0] n18452_o;
  wire [11:0] n18453_o;
  wire [31:0] alu_2_i_n18454;
  wire alu_2_i_n18455;
  wire [11:0] alu_2_i_n18456;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n18463_o;
  wire [11:0] n18464_o;
  wire [11:0] n18465_o;
  wire [31:0] alu_3_i_n18466;
  wire alu_3_i_n18467;
  wire [11:0] alu_3_i_n18468;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n18475_o;
  wire [11:0] n18476_o;
  wire [11:0] n18477_o;
  wire [31:0] alu_4_i_n18478;
  wire alu_4_i_n18479;
  wire [11:0] alu_4_i_n18480;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n18487_o;
  wire [11:0] n18488_o;
  wire [11:0] n18489_o;
  wire [31:0] alu_5_i_n18490;
  wire alu_5_i_n18491;
  wire [11:0] alu_5_i_n18492;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n18499_o;
  wire [11:0] n18500_o;
  wire [11:0] n18501_o;
  wire [31:0] alu_6_i_n18502;
  wire alu_6_i_n18503;
  wire [11:0] alu_6_i_n18504;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n18511_o;
  wire [11:0] n18512_o;
  wire [11:0] n18513_o;
  wire [31:0] alu_7_i_n18514;
  wire alu_7_i_n18515;
  wire [11:0] alu_7_i_n18516;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n18523_o;
  wire n18524_o;
  wire [12:0] ialu_i_n18525;
  wire ialu_i_n18526;
  wire ialu_i_n18527;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n18536;
  wire [95:0] register_bank_i_n18537;
  wire [16:0] n18538_o;
  wire [16:0] n18539_o;
  wire [95:0] register_bank_i_n18540;
  wire register_bank_i_n18541;
  wire register_bank_i_n18542;
  wire [2:0] register_bank_i_n18543;
  wire [2:0] register_bank_i_n18544;
  wire [1:0] register_bank_i_n18545;
  wire [2:0] register_bank_i_n18546;
  wire [2:0] register_bank_i_n18547;
  wire register_bank_i_n18548;
  wire [1:0] register_bank_i_n18549;
  wire [1:0] register_bank_i_n18550;
  wire register_bank_i_n18551;
  wire [1:0] register_bank_i_n18552;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n18585;
  wire instr_decoder2_i_n18586;
  wire [3:0] instr_decoder2_i_n18587;
  wire instr_decoder2_i_n18588;
  wire instr_decoder2_i_n18589;
  wire instr_decoder2_i_n18590;
  wire instr_decoder2_i_n18591;
  wire [11:0] instr_decoder2_i_n18592;
  wire [11:0] instr_decoder2_i_n18593;
  wire [11:0] instr_decoder2_i_n18594;
  wire instr_decoder2_i_n18595;
  wire instr_decoder2_i_n18596;
  wire instr_decoder2_i_n18597;
  wire [7:0] instr_decoder2_i_n18598;
  wire instr_decoder2_i_n18599;
  wire [11:0] instr_decoder2_i_n18600;
  wire instr_decoder2_i_n18601;
  wire instr_decoder2_i_n18602;
  wire [3:0] instr_decoder2_i_n18603;
  wire [3:0] instr_decoder2_i_n18604;
  wire instr_decoder2_i_n18605;
  wire instr_decoder2_i_n18606;
  wire [2:0] instr_decoder2_i_n18607;
  wire [12:0] instr_decoder2_i_n18608;
  wire instr_decoder2_i_n18609;
  wire [4:0] instr_decoder2_i_n18610;
  wire [12:0] instr_decoder2_i_n18611;
  wire [12:0] instr_decoder2_i_n18612;
  wire [7:0] instr_decoder2_i_n18613;
  wire [7:0] instr_decoder2_i_n18614;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n18675;
  wire instr_dispatch2_i1_n18676;
  wire [11:0] instr_dispatch2_i1_n18677;
  wire [11:0] instr_dispatch2_i1_n18678;
  wire instr_dispatch2_i1_n18679;
  wire instr_dispatch2_i1_n18680;
  wire instr_dispatch2_i1_n18681;
  wire instr_dispatch2_i1_n18682;
  wire instr_dispatch2_i1_n18683;
  wire instr_dispatch2_i1_n18684;
  wire instr_dispatch2_i1_n18685;
  wire instr_dispatch2_i1_n18686;
  wire [11:0] instr_dispatch2_i1_n18687;
  wire [7:0] instr_dispatch2_i1_n18688;
  wire [95:0] instr_dispatch2_i1_n18689;
  wire [7:0] instr_dispatch2_i1_n18690;
  wire [95:0] instr_dispatch2_i1_n18691;
  wire [95:0] instr_dispatch2_i1_n18692;
  wire [11:0] instr_dispatch2_i1_n18693;
  wire [4:0] instr_dispatch2_i1_n18694;
  wire [3:0] instr_dispatch2_i1_n18695;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n18741_o;
  wire [95:0] n18742_o;
  wire [7:0] n18743_o;
  wire [95:0] n18744_o;
  reg [95:0] n18745_q;
  wire [95:0] n18746_o;
  reg [95:0] n18747_q;
  reg n18748_q;
  reg n18749_q;
  wire n18750_o;
  reg n18751_q;
  wire [1:0] n18752_o;
  reg [1:0] n18753_q;
  wire [1:0] n18754_o;
  reg [1:0] n18755_q;
  wire [2:0] n18756_o;
  reg [2:0] n18757_q;
  wire [2:0] n18758_o;
  reg [2:0] n18759_q;
  wire n18760_o;
  reg n18761_q;
  wire [1:0] n18762_o;
  reg [1:0] n18763_q;
  reg [2:0] n18764_q;
  reg [2:0] n18765_q;
  reg [1:0] n18766_q;
  reg [2:0] n18769_q;
  reg [2:0] n18770_q;
  reg n18771_q;
  reg [1:0] n18772_q;
  reg [1:0] n18773_q;
  reg n18774_q;
  reg [1:0] n18775_q;
  reg [21:0] n18776_q;
  reg [2:0] n18777_q;
  reg [21:0] n18778_q;
  reg [95:0] n18779_q;
  wire n18780_o;
  reg n18781_q;
  wire n18782_o;
  reg n18783_q;
  wire n18784_o;
  reg n18785_q;
  reg [21:0] n18788_q;
  reg [21:0] n18789_q;
  wire [5:0] n18790_o;
  reg [5:0] n18791_q;
  wire n18792_o;
  reg n18793_q;
  wire [2:0] n18796_o;
  reg [2:0] n18797_q;
  wire [1:0] n18798_o;
  reg [1:0] n18799_q;
  wire n18800_o;
  reg n18801_q;
  wire [21:0] n18802_o;
  reg [21:0] n18803_q;
  wire n18804_o;
  reg n18805_q;
  wire [2:0] n18806_o;
  reg [2:0] n18807_q;
  wire [1:0] n18808_o;
  reg [1:0] n18809_q;
  wire n18810_o;
  wire n18811_o;
  wire n18812_o;
  reg n18813_q;
  wire n18814_o;
  wire n18815_o;
  wire [21:0] n18816_o;
  reg [21:0] n18817_q;
  wire n18818_o;
  reg n18819_q;
  wire [1:0] n18820_o;
  reg [1:0] n18821_q;
  wire [1:0] n18822_o;
  reg [1:0] n18823_q;
  wire n18824_o;
  reg n18825_q;
  wire [1:0] n18826_o;
  reg [1:0] n18827_q;
  reg [83:0] n18828_q;
  wire [95:0] n18829_o;
  reg [2:0] n18830_q;
  reg [2:0] n18831_q;
  reg [2:0] n18832_q;
  reg [79:0] n18834_q;
  reg [31:0] n18835_q;
  reg n18836_q;
  reg n18837_q;
  reg n18838_q;
  reg [1:0] n18839_q;
  reg [3:0] n18840_q;
  reg n18841_q;
  reg [3:0] n18842_q;
  reg n18843_q;
  reg [3:0] n18844_q;
  reg n18845_q;
  reg n18846_q;
  reg [1:0] n18847_q;
  reg [27:0] n18848_q;
  reg n18849_q;
  reg n18850_q;
  reg n18852_q;
  reg n18853_q;
  reg n18855_q;
  reg n18856_q;
  reg n18857_q;
  reg [21:0] n18858_q;
  reg n18859_q;
  reg [21:0] n18860_q;
  reg [21:0] n18861_q;
  reg n18862_q;
  reg [21:0] n18863_q;
  reg [5:0] n18864_q;
  reg n18865_q;
  reg n18866_q;
  reg n18867_q;
  reg [2:0] n18868_q;
  reg [1:0] n18869_q;
  reg n18870_q;
  reg n18871_q;
  reg [2:0] n18872_q;
  reg [1:0] n18873_q;
  reg n18874_q;
  reg [1:0] n18875_q;
  reg [1:0] n18876_q;
  reg n18877_q;
  reg [1:0] n18878_q;
  reg [95:0] n18879_q;
  reg n18880_q;
  wire [2:0] n18881_o;
  wire [2:0] n18882_o;
  assign i_y_neg_out = n18523_o;
  assign i_y_zero_out = n18524_o;
  assign dp_readdata_out = n18196_o;
  assign dp_readdata_vm_out = n18198_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n18881_o;
  assign dp_read_vaddr_out = n18882_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n18176_o;
  assign dp_read_data_type_out = n18178_o;
  assign dp_read_stream_out = n18180_o;
  assign dp_read_stream_id_out = n18182_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n18536; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n18537; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n18675; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n18676; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n18684; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n18681; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n18682; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n18683; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n18689; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n18690; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n18592; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n18593; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n18594; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n18374; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n18609; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n18585; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n18691; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n18692; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n18693; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n18741_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n18742_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n18743_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n18694; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n18695; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n18587; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n18424_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n18397_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n18190_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n18677; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n18678; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n18687; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n18688; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n18188_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n18189_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n18586; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n18591; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n18588; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n18589; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n18590; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n18599; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n18600; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n18595; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n18596; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n18597; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n18598; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n18679; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n18680; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n18686; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n18601; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n18602; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n18603; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n18373; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n18604; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n18605; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n18606; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n18607; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n18608; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n18745_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n18747_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n18748_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n18749_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n18751_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n18753_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n18755_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n18757_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n18759_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n18761_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n18763_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n18610; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n18611; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n18612; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n18525; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n18526; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n18527; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n18685; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n18613; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n18614; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n18367; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n18368; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n17856_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n17857_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n17896_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n17858_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n17898_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n17899_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n17900_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n17901_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n17902_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n17903_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n17904_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n17859_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n17860_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n17861_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n17862_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n17863_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n17864_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n17865_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n17866_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n17867_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n17868_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n18150_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n17869_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n17870_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n17906_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n17909_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n18764_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n18765_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n18766_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n18769_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n18770_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n18771_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n18772_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n18773_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n18774_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n18775_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n18776_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n18777_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n18778_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n18779_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n18781_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n18783_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n18785_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n18788_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n18789_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n18791_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n18793_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n18797_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n18799_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n18801_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n18803_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n18805_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n18807_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n18809_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n18813_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n18817_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n18819_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n18821_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n18823_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n18825_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n18827_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n18829_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n18830_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n18831_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n18832_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n18174_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n17835_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n18542; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n18543; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n18544; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n18545; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n18546; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n18547; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n18540; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n18541; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n18548; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n18549; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n18550; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n18551; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n18552; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n17713_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n17714_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n17715_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n18834_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n18835_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n18836_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n18837_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n18838_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n18839_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n18840_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n18841_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n18842_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n18843_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n18844_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n18845_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n18846_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n18847_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n18848_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n18849_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n18850_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n18852_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n18853_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n18855_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n18856_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n18857_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n18858_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n18859_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n18860_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n18861_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n18862_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n18863_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n18864_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n18865_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n18866_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n18867_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n18868_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n18869_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n18870_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n18871_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n18872_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n18873_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n18874_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n18875_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n18876_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n18877_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n18878_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n18879_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n18880_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n17713_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n17714_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n17715_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n17718_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n17806_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n17807_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n17808_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n17809_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n17812_o = n17809_o ? 3'b000 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n17814_o = n17808_o + n17806_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n17815_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n17816_o = n17815_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n17817_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n17818_o = n17817_o & n17816_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n17819_o = n17806_o & n17808_o;
  /* ../../HW/src/pcore/pcore.vhd:215:8  */
  assign n17820_o = {n17812_o, 2'b01};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n17821_o = n17806_o & n17820_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n17822_o = n17819_o == n17821_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n17823_o = n17822_o & n17807_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n17824_o = ~n17807_o;
  /* ../../HW/src/pcore/pcore.vhd:106:8  */
  assign n17825_o = {n17812_o, 2'b01};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n17826_o = $unsigned(n17825_o) >= $unsigned(n17808_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n17827_o = n17826_o & n17824_o;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n17828_o = {n17812_o, 2'b01};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n17829_o = $unsigned(n17828_o) <= $unsigned(n17814_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n17830_o = n17829_o & n17827_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n17831_o = n17823_o | n17830_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n17832_o = n17831_o & n17818_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n17835_o = n17832_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n17841_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n17843_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n17845_o = n17843_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n17847_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n17848_o = n17847_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n17849_o = dp_read_gen_valid_in_r & n17848_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n17851_o = n17849_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n17853_o = n17849_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n17855_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17856_o = n17841_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17857_o = n17841_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17858_o = n17841_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17859_o = n17841_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17860_o = n17841_o ? n17845_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17861_o = n17841_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17862_o = n17841_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17863_o = n17841_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17864_o = n17841_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17865_o = n17841_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17866_o = n17841_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17867_o = n17841_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17868_o = n17841_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17869_o = n17841_o ? n17851_o : n17855_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n17870_o = n17841_o ? n17853_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n17875_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n17876_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n17877_o = dp_write_in_r & n17876_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n17878_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n17879_o = n17877_o & n17878_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n17881_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n17883_o = n17881_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n17885_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n17886_o = n17885_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n17887_o = dp_write_gen_valid_in_r & n17886_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n17889_o = n17887_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n17893_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n17895_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17896_o = n17875_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17898_o = n17875_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17899_o = n17875_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17900_o = n17875_o ? n17879_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17901_o = n17875_o ? n17883_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17902_o = n17875_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17903_o = n17875_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17904_o = n17875_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17906_o = n17875_o ? n17889_o : n17893_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n17909_o = n17875_o ? 3'b000 : n17895_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n17914_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n17917_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n17918_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n17919_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n17921_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n17922_o = n17918_o ? n17919_o : n17921_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n17924_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n17925_o = n17917_o ? n17922_o : n17924_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n17927_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n17991_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n18060_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n18063_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n18064_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n18065_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n18067_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n18068_o = n18064_o ? n18065_o : n18067_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n18070_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n18071_o = n18063_o ? n18068_o : n18070_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n18073_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n18074_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n18075_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n18085_o = n18073_o ? n18074_o : n18075_o;
  assign n18127_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n18128_o = n18060_o ? 12'b000000000000 : n18127_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n18142_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n18144_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n18145_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n18146_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n18147_o = n18144_o ? n18145_o : n18146_o;
  assign n18149_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n18147_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n18150_o = n18142_o ? n18149_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n18156_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n18157_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n18158_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n18160_o = n18156_o == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n18161_o = n18160_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n18163_o = n18157_o == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n18164_o = n18163_o & n18161_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n18167_o = n18164_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n18169_o = n18156_o == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n18170_o = n18169_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n18173_o = n18170_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n18174_o = n18158_o ? n18167_o : n18173_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n18176_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n18178_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n18180_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n18182_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n18188_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n18189_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n18190_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n18193_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n18194_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n18196_o = n18193_o ? 96'bZ : n18194_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n18198_o = n18193_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n18203_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n18254_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n18257_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n18258_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n18259_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n18261_o = n18258_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n18262_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n18264_o = n18258_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n18265_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n18267_o = n18258_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n18268_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n18270_o = n18258_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n18271_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n18273_o = n18258_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n18274_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n18276_o = n18258_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n18277_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n18279_o = n18258_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n18280_o = dp_readdata_vm[11:0];
  assign n18281_o = {n18279_o, n18276_o, n18273_o, n18270_o, n18267_o, n18264_o, n18261_o};
  assign n18282_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18283_o = n18282_o;
      7'b0100000: n18283_o = n18282_o;
      7'b0010000: n18283_o = n18282_o;
      7'b0001000: n18283_o = n18282_o;
      7'b0000100: n18283_o = n18282_o;
      7'b0000010: n18283_o = n18282_o;
      7'b0000001: n18283_o = n18282_o;
      default: n18283_o = n18280_o;
    endcase
  assign n18284_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18285_o = n18277_o;
      7'b0100000: n18285_o = n18284_o;
      7'b0010000: n18285_o = n18284_o;
      7'b0001000: n18285_o = n18284_o;
      7'b0000100: n18285_o = n18284_o;
      7'b0000010: n18285_o = n18284_o;
      7'b0000001: n18285_o = n18284_o;
      default: n18285_o = n18284_o;
    endcase
  assign n18286_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18287_o = n18286_o;
      7'b0100000: n18287_o = n18274_o;
      7'b0010000: n18287_o = n18286_o;
      7'b0001000: n18287_o = n18286_o;
      7'b0000100: n18287_o = n18286_o;
      7'b0000010: n18287_o = n18286_o;
      7'b0000001: n18287_o = n18286_o;
      default: n18287_o = n18286_o;
    endcase
  assign n18288_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18289_o = n18288_o;
      7'b0100000: n18289_o = n18288_o;
      7'b0010000: n18289_o = n18271_o;
      7'b0001000: n18289_o = n18288_o;
      7'b0000100: n18289_o = n18288_o;
      7'b0000010: n18289_o = n18288_o;
      7'b0000001: n18289_o = n18288_o;
      default: n18289_o = n18288_o;
    endcase
  assign n18290_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18291_o = n18290_o;
      7'b0100000: n18291_o = n18290_o;
      7'b0010000: n18291_o = n18290_o;
      7'b0001000: n18291_o = n18268_o;
      7'b0000100: n18291_o = n18290_o;
      7'b0000010: n18291_o = n18290_o;
      7'b0000001: n18291_o = n18290_o;
      default: n18291_o = n18290_o;
    endcase
  assign n18292_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18293_o = n18292_o;
      7'b0100000: n18293_o = n18292_o;
      7'b0010000: n18293_o = n18292_o;
      7'b0001000: n18293_o = n18292_o;
      7'b0000100: n18293_o = n18265_o;
      7'b0000010: n18293_o = n18292_o;
      7'b0000001: n18293_o = n18292_o;
      default: n18293_o = n18292_o;
    endcase
  assign n18294_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18295_o = n18294_o;
      7'b0100000: n18295_o = n18294_o;
      7'b0010000: n18295_o = n18294_o;
      7'b0001000: n18295_o = n18294_o;
      7'b0000100: n18295_o = n18294_o;
      7'b0000010: n18295_o = n18262_o;
      7'b0000001: n18295_o = n18294_o;
      default: n18295_o = n18294_o;
    endcase
  assign n18296_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n18281_o)
      7'b1000000: n18297_o = n18296_o;
      7'b0100000: n18297_o = n18296_o;
      7'b0010000: n18297_o = n18296_o;
      7'b0001000: n18297_o = n18296_o;
      7'b0000100: n18297_o = n18296_o;
      7'b0000010: n18297_o = n18296_o;
      7'b0000001: n18297_o = n18259_o;
      default: n18297_o = n18296_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n18299_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n18302_o = n18299_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n18303_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n18304_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n18305_o = {n18297_o, n18295_o, n18293_o, n18291_o, n18289_o, n18287_o, n18285_o, n18283_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n18306_o = n18257_o ? n18305_o : n18303_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n18307_o = n18257_o ? dp_readdata2_r : n18304_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n18309_o = n18257_o ? n18302_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n18311_o = n18257_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n18313_o = n18257_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n18318_o = dp_readena_vm ? n18309_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n18367 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n18368 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n18373 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n18374 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n18381_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n18383_o = dp_rd_pid == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n18384_o = n18383_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n18386_o = dp_rd_cid == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n18387_o = n18386_o & n18384_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n18390_o = n18387_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n18392_o = dp_rd_pid == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n18393_o = n18392_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n18396_o = n18393_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n18397_o = n18381_o ? n18390_o : n18396_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n18405_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n18406_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n18407_o = dp_mcast_addr + n18405_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n18408_o = n18405_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n18410_o = n18405_o & 5'b00001;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n18411_o = n18408_o == n18410_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n18412_o = n18411_o & n18406_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n18413_o = ~n18406_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n18415_o = $unsigned(5'b00001) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n18416_o = n18415_o & n18413_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n18418_o = $unsigned(5'b00001) <= $unsigned(n18407_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n18419_o = n18418_o & n18416_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n18420_o = n18412_o | n18419_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n18421_o = n18420_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n18424_o = n18421_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n18427_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n18428_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n18429_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n18430 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n18431 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n18432 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18427_o),
    .x1_in(n18428_o),
    .x2_in(n18429_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n18439_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n18440_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n18441_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n18442 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n18443 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n18444 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18439_o),
    .x1_in(n18440_o),
    .x2_in(n18441_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n18451_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n18452_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n18453_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n18454 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n18455 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n18456 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18451_o),
    .x1_in(n18452_o),
    .x2_in(n18453_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n18463_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n18464_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n18465_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n18466 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n18467 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n18468 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18463_o),
    .x1_in(n18464_o),
    .x2_in(n18465_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n18475_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n18476_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n18477_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n18478 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n18479 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n18480 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18475_o),
    .x1_in(n18476_o),
    .x2_in(n18477_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n18487_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n18488_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n18489_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n18490 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n18491 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n18492 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18487_o),
    .x1_in(n18488_o),
    .x2_in(n18489_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n18499_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n18500_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n18501_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n18502 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n18503 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n18504 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18499_o),
    .x1_in(n18500_o),
    .x2_in(n18501_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n18511_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n18512_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n18513_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n18514 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n18515 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n18516 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n18511_o),
    .x1_in(n18512_o),
    .x2_in(n18513_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n18523_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n18524_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n18525 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n18526 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n18527 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n18536 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n18537 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n18538_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n18539_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n18540 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n18541 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n18542 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n18543 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n18544 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n18545 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n18546 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n18547 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n18548 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n18549 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n18550 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n18551 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n18552 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n18538_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n18539_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n18585 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n18586 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n18587 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n18588 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n18589 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n18590 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n18591 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n18592 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n18593 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n18594 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n18595 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n18596 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n18597 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n18598 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n18599 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n18600 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n18601 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n18602 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n18603 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n18604 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n18605 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n18606 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n18607 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n18608 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n18609 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n18610 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n18611 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n18612 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n18613 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n18614 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_0_1 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n18675 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n18676 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n18677 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n18678 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n18679 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n18680 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n18681 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n18682 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n18683 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n18684 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n18685 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n18686 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n18687 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n18688 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n18689 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n18690 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n18691 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n18692 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n18693 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n18694 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n18695 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n18741_o = {alu_7_i_n18514, alu_6_i_n18502, alu_5_i_n18490, alu_4_i_n18478, alu_3_i_n18466, alu_2_i_n18454, alu_1_i_n18442, alu_0_i_n18430};
  assign n18742_o = {alu_7_i_n18516, alu_6_i_n18504, alu_5_i_n18492, alu_4_i_n18480, alu_3_i_n18468, alu_2_i_n18456, alu_1_i_n18444, alu_0_i_n18432};
  assign n18743_o = {alu_7_i_n18515, alu_6_i_n18503, alu_5_i_n18491, alu_4_i_n18479, alu_3_i_n18467, alu_2_i_n18455, alu_1_i_n18443, alu_0_i_n18431};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18744_o = dp_readena_vm ? n18306_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18745_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n18745_q <= n18744_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18746_o = dp_readena_vm ? n18307_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18747_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n18747_q <= n18746_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18748_q <= 1'b0;
    else
      n18748_q <= n18318_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18749_q <= 1'b0;
    else
      n18749_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18750_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18751_q <= 1'b0;
    else
      n18751_q <= n18750_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18752_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18753_q <= 2'b00;
    else
      n18753_q <= n18752_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18754_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18755_q <= 2'b00;
    else
      n18755_q <= n18754_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18756_o = dp_readena_vm ? n18311_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18757_q <= 3'b000;
    else
      n18757_q <= n18756_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18758_o = dp_readena_vm ? n18313_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18759_q <= 3'b000;
    else
      n18759_q <= n18758_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18760_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18761_q <= 1'b0;
    else
      n18761_q <= n18760_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n18762_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n18254_o)
    if (n18254_o)
      n18763_q <= 2'b00;
    else
      n18763_q <= n18762_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18764_q <= 3'b000;
    else
      n18764_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18765_q <= 3'b000;
    else
      n18765_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18766_q <= 2'b00;
    else
      n18766_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18769_q <= 3'b000;
    else
      n18769_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18770_q <= 3'b000;
    else
      n18770_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18771_q <= 1'b0;
    else
      n18771_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18772_q <= 2'b00;
    else
      n18772_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18773_q <= 2'b00;
    else
      n18773_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18774_q <= 1'b0;
    else
      n18774_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18775_q <= 2'b00;
    else
      n18775_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18776_q <= 22'b0000000000000000000000;
    else
      n18776_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18777_q <= 3'b000;
    else
      n18777_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18778_q <= 22'b0000000000000000000000;
    else
      n18778_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18779_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n18779_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18780_o = n17927_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18781_q <= 1'b0;
    else
      n18781_q <= n18780_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18782_o = n17927_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18783_q <= 1'b0;
    else
      n18783_q <= n18782_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18784_o = n18073_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18785_q <= 1'b0;
    else
      n18785_q <= n18784_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18788_q <= 22'b0000000000000000000000;
    else
      n18788_q <= n17925_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18789_q <= 22'b0000000000000000000000;
    else
      n18789_q <= n18071_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18790_o = n18073_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18791_q <= 6'b000000;
    else
      n18791_q <= n18790_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18792_o = n18073_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18793_q <= 1'b0;
    else
      n18793_q <= n18792_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18796_o = n18073_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18797_q <= 3'b000;
    else
      n18797_q <= n18796_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18798_o = n18073_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18799_q <= 2'b00;
    else
      n18799_q <= n18798_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18800_o = n18073_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18801_q <= 1'b0;
    else
      n18801_q <= n18800_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n18802_o = n18073_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18803_q <= 22'b0000000000000000000000;
    else
      n18803_q <= n18802_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18804_o = n17927_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18805_q <= 1'b0;
    else
      n18805_q <= n18804_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18806_o = n17927_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18807_q <= 3'b000;
    else
      n18807_q <= n18806_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18808_o = n17927_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18809_q <= 2'b00;
    else
      n18809_q <= n18808_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n18810_o = ~n17914_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n18811_o = n17927_o & n18810_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18812_o = n18811_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n18813_q <= n18812_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n18814_o = ~n17914_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n18815_o = n17927_o & n18814_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18816_o = n18815_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n18817_q <= n18816_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18818_o = n17927_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18819_q <= 1'b0;
    else
      n18819_q <= n18818_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18820_o = n17927_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18821_q <= 2'b00;
    else
      n18821_q <= n18820_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18822_o = n17927_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18823_q <= 2'b00;
    else
      n18823_q <= n18822_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18824_o = n17927_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18825_q <= 1'b0;
    else
      n18825_q <= n18824_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n18826_o = n17927_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18827_q <= 2'b00;
    else
      n18827_q <= n18826_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18828_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n18828_q <= n18085_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n18829_o = {n18128_o, n18828_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18830_q <= 3'b000;
    else
      n18830_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n17914_o)
    if (n17914_o)
      n18831_q <= 3'b000;
    else
      n18831_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n18060_o)
    if (n18060_o)
      n18832_q <= 3'b000;
    else
      n18832_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18834_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n18834_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18835_q <= 32'b00000000000000000000000000000000;
    else
      n18835_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18836_q <= 1'b0;
    else
      n18836_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18837_q <= 1'b0;
    else
      n18837_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18838_q <= 1'b0;
    else
      n18838_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18839_q <= 2'b00;
    else
      n18839_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18840_q <= 4'b0000;
    else
      n18840_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18841_q <= 1'b0;
    else
      n18841_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18842_q <= 4'b0000;
    else
      n18842_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18843_q <= 1'b0;
    else
      n18843_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18844_q <= 4'b0000;
    else
      n18844_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18845_q <= 1'b0;
    else
      n18845_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18846_q <= 1'b0;
    else
      n18846_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18847_q <= 2'b00;
    else
      n18847_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n18203_o)
    if (n18203_o)
      n18848_q <= 28'b0000000000000000000000000000;
    else
      n18848_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18849_q <= 1'b0;
    else
      n18849_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18850_q <= 1'b0;
    else
      n18850_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18852_q <= 1'b0;
    else
      n18852_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n17991_o)
    if (n17991_o)
      n18853_q <= 1'b0;
    else
      n18853_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18855_q <= 1'b0;
    else
      n18855_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18856_q <= 1'b0;
    else
      n18856_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18857_q <= 1'b0;
    else
      n18857_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18858_q <= 22'b0000000000000000000000;
    else
      n18858_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18859_q <= 1'b0;
    else
      n18859_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18860_q <= 22'b0000000000000000000000;
    else
      n18860_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18861_q <= 22'b0000000000000000000000;
    else
      n18861_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18862_q <= 1'b0;
    else
      n18862_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18863_q <= 22'b0000000000000000000000;
    else
      n18863_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18864_q <= 6'b000000;
    else
      n18864_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18865_q <= 1'b0;
    else
      n18865_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18866_q <= 1'b0;
    else
      n18866_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18867_q <= 1'b0;
    else
      n18867_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18868_q <= 3'b000;
    else
      n18868_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18869_q <= 2'b00;
    else
      n18869_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18870_q <= 1'b0;
    else
      n18870_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18871_q <= 1'b0;
    else
      n18871_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18872_q <= 3'b000;
    else
      n18872_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18873_q <= 2'b00;
    else
      n18873_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18874_q <= 1'b0;
    else
      n18874_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18875_q <= 2'b00;
    else
      n18875_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18876_q <= 2'b00;
    else
      n18876_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18877_q <= 1'b0;
    else
      n18877_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18878_q <= 2'b00;
    else
      n18878_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18879_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n18879_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n17718_o)
    if (n17718_o)
      n18880_q <= 1'b0;
    else
      n18880_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n18881_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n18882_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module pcore_0_0
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_share_in,
   input  dp_rd_fork_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in_in,
   output i_y_neg_out,
   output i_y_zero_out,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output dp_readena_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out);
  wire [95:0] rd_x1_data1;
  wire [95:0] rd_x2_data1;
  wire rd_en1;
  wire rd_vm;
  wire wr_en1;
  wire wr_xreg1;
  wire wr_flag1;
  wire wr_xreg_flag1;
  wire [95:0] wr_data1;
  wire [7:0] wr_vector_lane;
  wire [11:0] x1_addr1;
  wire [11:0] x2_addr1;
  wire [11:0] y_addr1;
  wire [12:0] rd_lane;
  wire wr_lane;
  wire [4:0] opcode1;
  wire [95:0] mu_x1;
  wire [95:0] mu_x2;
  wire [11:0] mu_x_scalar;
  wire [255:0] mu_y;
  wire [95:0] mu_y2;
  wire [7:0] mu_result;
  wire [4:0] mu_opcodes;
  wire [3:0] mu_tid;
  wire [3:0] tid_decoder2dispatch;
  wire write;
  wire read;
  wire [4:0] dp_mcast_addr;
  wire [11:0] rd_x1_addr1;
  wire [11:0] rd_x2_addr1;
  wire [11:0] wr_addr1;
  wire [7:0] wr_result_addr1;
  wire [1:0] dp_rd_pid;
  wire [2:0] dp_rd_cid;
  wire en1;
  wire mu_vm;
  wire mu_xreg1;
  wire mu_flag1;
  wire mu_wren;
  wire x1_c1_en;
  wire [11:0] x1_c1;
  wire x1_vector;
  wire x2_vector;
  wire y_vector;
  wire [7:0] vector_lane;
  wire rd_x1_vector1;
  wire rd_x2_vector1;
  wire wr_vector;
  wire i_rd_en1;
  wire i_rd_vm;
  wire [3:0] i_rd_tid1;
  wire [103:0] i_rd_data1;
  wire [3:0] i_wr_tid1;
  wire i_wr_en1;
  wire i_wr_vm;
  wire [2:0] i_wr_addr1;
  wire [12:0] i_wr_data1;
  wire [95:0] dp_readdata_r;
  wire [95:0] dp_readdata2_r;
  wire dp_readena_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid2_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_type2_r;
  wire [2:0] dp_read_vector2_r;
  wire [2:0] dp_read_vaddr2_r;
  wire dp_read_stream2_r;
  wire [1:0] dp_read_stream_id2_r;
  wire [4:0] i_opcode;
  wire [12:0] i_x1;
  wire [12:0] i_x2;
  wire [12:0] i_y;
  wire i_y_neg;
  wire i_y_zero;
  wire wr_vm;
  wire [7:0] result_write_addr;
  wire [7:0] result_raddr1;
  wire [7:0] result_waddr1;
  wire [12:0] result_read;
  wire [255:0] xreg_read;
  wire dp_rd_vm;
  wire dp_rd_fork;
  wire dp_wr_vm;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_wr_addr;
  wire [5:0] dp_wr_mcast;
  wire dp_write;
  wire [2:0] dp_write_vector;
  wire [1:0] dp_write_scatter;
  wire dp_write_share;
  wire [21:0] dp_write_step;
  wire dp_read;
  wire [2:0] dp_read_vector;
  wire [1:0] dp_read_scatter;
  wire dp_read_share;
  wire [21:0] dp_read_step;
  wire dp_read_gen_valid;
  wire [1:0] dp_read_data_flow;
  wire [1:0] dp_read_data_type;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_writedata;
  wire [2:0] read_scatter_cnt;
  wire [2:0] read_scatter_vector;
  wire [2:0] write_scatter_cnt;
  wire [2:0] write_scatter_curr;
  wire [2:0] write_scatter_curr_r;
  wire [2:0] gen_read_vector_r;
  wire [1:0] gen_read_scatter_r;
  wire [2:0] gen_read_scatter_cnt_r;
  wire [2:0] gen_read_scatter_vector_r;
  wire gen_read_gen_valid_r;
  wire [1:0] gen_read_data_flow_r;
  wire [1:0] gen_read_data_type_r;
  wire gen_read_stream_r;
  wire [1:0] gen_read_stream_id_r;
  wire [21:0] gen_rd_addr_r;
  wire [2:0] gen_write_vector_r;
  wire [21:0] gen_wr_addr_r;
  wire [95:0] gen_writedata_r;
  wire dp_rd_vm_r;
  wire dp_rd_fork_r;
  wire dp_wr_vm_r;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_wr_addr_r;
  wire [5:0] dp_wr_mcast_r;
  wire dp_write_r;
  wire [2:0] dp_write_vector_r;
  wire [1:0] dp_write_scatter_r;
  wire dp_write_share_r;
  wire [21:0] dp_write_step_r;
  wire dp_read_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire dp_read_share_r;
  wire [21:0] dp_read_step_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [95:0] dp_writedata_r;
  wire [2:0] read_scatter_cnt_r;
  wire [2:0] read_scatter_vector_r;
  wire [2:0] write_scatter_cnt_r;
  wire read_match;
  wire write_match;
  wire dp_readena_vm;
  wire [2:0] dp_read_vector_vm;
  wire [2:0] dp_read_vaddr_vm;
  wire [1:0] dp_read_scatter_vm;
  wire [2:0] dp_read_scatter_cnt_vm;
  wire [2:0] dp_read_scatter_vector_vm;
  wire [95:0] dp_readdata_vm;
  wire dp_readdata_vm_vm;
  wire dp_read_gen_valid_vm;
  wire [1:0] dp_read_data_flow_vm;
  wire [1:0] dp_read_data_type_vm;
  wire dp_read_stream_vm;
  wire [1:0] dp_read_stream_id_vm;
  wire tid_valid1;
  wire pre_tid_valid1;
  wire pre_pre_tid_valid1;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire vm_r;
  wire [1:0] data_model_r;
  wire [3:0] tid_r;
  wire tid_valid1_r;
  wire [3:0] pre_tid_r;
  wire pre_tid_valid1_r;
  wire [3:0] pre_pre_tid_r;
  wire pre_pre_tid_valid1_r;
  wire pre_pre_vm_r;
  wire [1:0] pre_pre_data_model_r;
  wire [27:0] pre_iregister_auto_r;
  wire gen_write_r;
  wire gen_write_vm_r;
  wire gen_read_r;
  wire gen_read_vm_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_rd_step_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_wr_share_in_r;
  wire [21:0] dp_wr_step_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_wr_fork_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_rd_fork_in_r;
  wire dp_read_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n16531_o;
  wire n16532_o;
  wire n16533_o;
  wire n16536_o;
  wire [4:0] n16624_o;
  wire n16625_o;
  wire [4:0] n16626_o;
  wire n16627_o;
  wire [2:0] n16630_o;
  wire [4:0] n16632_o;
  wire n16633_o;
  wire n16634_o;
  wire n16635_o;
  wire n16636_o;
  wire [4:0] n16637_o;
  wire [4:0] n16638_o;
  wire [4:0] n16639_o;
  wire n16640_o;
  wire n16641_o;
  wire n16642_o;
  wire [4:0] n16643_o;
  wire n16644_o;
  wire n16645_o;
  wire [4:0] n16646_o;
  wire n16647_o;
  wire n16648_o;
  wire n16649_o;
  wire n16650_o;
  wire n16653_o;
  wire n16659_o;
  wire n16661_o;
  wire [2:0] n16663_o;
  wire n16665_o;
  wire n16666_o;
  wire n16667_o;
  wire [2:0] n16669_o;
  wire [2:0] n16671_o;
  wire [2:0] n16673_o;
  wire n16674_o;
  wire n16675_o;
  wire [21:0] n16676_o;
  wire n16677_o;
  wire [2:0] n16678_o;
  wire [1:0] n16679_o;
  wire n16680_o;
  wire [21:0] n16681_o;
  wire n16682_o;
  wire [1:0] n16683_o;
  wire [1:0] n16684_o;
  wire n16685_o;
  wire [1:0] n16686_o;
  wire [2:0] n16687_o;
  wire [2:0] n16688_o;
  wire n16693_o;
  wire n16694_o;
  wire n16695_o;
  wire n16696_o;
  wire n16697_o;
  wire n16699_o;
  wire [2:0] n16701_o;
  wire n16703_o;
  wire n16704_o;
  wire n16705_o;
  wire [2:0] n16707_o;
  wire [2:0] n16711_o;
  wire [2:0] n16713_o;
  wire n16714_o;
  wire [21:0] n16716_o;
  wire [5:0] n16717_o;
  wire n16718_o;
  wire [2:0] n16719_o;
  wire [1:0] n16720_o;
  wire n16721_o;
  wire [21:0] n16722_o;
  wire [2:0] n16724_o;
  wire [2:0] n16727_o;
  wire n16732_o;
  wire n16735_o;
  wire n16736_o;
  wire [21:0] n16737_o;
  wire [21:0] n16739_o;
  wire [21:0] n16740_o;
  wire [21:0] n16742_o;
  wire [21:0] n16743_o;
  wire n16745_o;
  wire n16809_o;
  wire n16878_o;
  wire n16881_o;
  wire n16882_o;
  wire [21:0] n16883_o;
  wire [21:0] n16885_o;
  wire [21:0] n16886_o;
  wire [21:0] n16888_o;
  wire [21:0] n16889_o;
  wire n16891_o;
  wire [83:0] n16892_o;
  wire [83:0] n16893_o;
  wire [83:0] n16903_o;
  wire [11:0] n16945_o;
  wire [11:0] n16946_o;
  wire n16960_o;
  wire n16962_o;
  wire [11:0] n16963_o;
  wire [11:0] n16964_o;
  wire [11:0] n16965_o;
  wire [95:0] n16967_o;
  wire [95:0] n16968_o;
  wire [1:0] n16974_o;
  wire [2:0] n16975_o;
  wire n16976_o;
  wire n16978_o;
  wire n16979_o;
  wire n16981_o;
  wire n16982_o;
  wire n16985_o;
  wire n16987_o;
  wire n16988_o;
  wire n16991_o;
  wire n16992_o;
  wire [1:0] n16994_o;
  wire [1:0] n16996_o;
  wire n16998_o;
  wire [1:0] n17000_o;
  wire [1:0] n17006_o;
  wire [2:0] n17007_o;
  wire [4:0] n17008_o;
  wire n17011_o;
  wire [95:0] n17012_o;
  wire [95:0] n17014_o;
  wire n17016_o;
  wire n17021_o;
  wire n17072_o;
  wire n17075_o;
  wire [2:0] n17076_o;
  wire [11:0] n17077_o;
  wire n17079_o;
  wire [11:0] n17080_o;
  wire n17082_o;
  wire [11:0] n17083_o;
  wire n17085_o;
  wire [11:0] n17086_o;
  wire n17088_o;
  wire [11:0] n17089_o;
  wire n17091_o;
  wire [11:0] n17092_o;
  wire n17094_o;
  wire [11:0] n17095_o;
  wire n17097_o;
  wire [11:0] n17098_o;
  wire [6:0] n17099_o;
  wire [11:0] n17100_o;
  reg [11:0] n17101_o;
  wire [11:0] n17102_o;
  reg [11:0] n17103_o;
  wire [11:0] n17104_o;
  reg [11:0] n17105_o;
  wire [11:0] n17106_o;
  reg [11:0] n17107_o;
  wire [11:0] n17108_o;
  reg [11:0] n17109_o;
  wire [11:0] n17110_o;
  reg [11:0] n17111_o;
  wire [11:0] n17112_o;
  reg [11:0] n17113_o;
  wire [11:0] n17114_o;
  reg [11:0] n17115_o;
  wire n17117_o;
  wire n17120_o;
  wire [95:0] n17121_o;
  wire [95:0] n17122_o;
  wire [95:0] n17123_o;
  wire [95:0] n17124_o;
  wire [95:0] n17125_o;
  wire n17127_o;
  wire [2:0] n17129_o;
  wire [2:0] n17131_o;
  wire n17136_o;
  wire [12:0] xregister_file_i_n17185;
  wire [255:0] xregister_file_i_n17186;
  wire [12:0] xregister_file_i_read_result_out;
  wire [255:0] xregister_file_i_read_xreg_out;
  wire [103:0] iregister_i_n17191;
  wire [12:0] iregister_i_n17192;
  wire [103:0] iregister_i_rd_data1_out;
  wire [12:0] iregister_i_rd_lane_out;
  wire n17199_o;
  wire n17201_o;
  wire n17202_o;
  wire n17204_o;
  wire n17205_o;
  wire n17208_o;
  wire n17210_o;
  wire n17211_o;
  wire n17214_o;
  wire n17215_o;
  wire [4:0] n17223_o;
  wire n17224_o;
  wire [4:0] n17225_o;
  wire [4:0] n17226_o;
  wire [4:0] n17228_o;
  wire n17229_o;
  wire n17230_o;
  wire n17231_o;
  wire n17233_o;
  wire n17234_o;
  wire n17236_o;
  wire n17237_o;
  wire n17238_o;
  wire n17239_o;
  wire n17242_o;
  wire [31:0] n17245_o;
  wire [11:0] n17246_o;
  wire [11:0] n17247_o;
  wire [31:0] alu_0_i_n17248;
  wire alu_0_i_n17249;
  wire [11:0] alu_0_i_n17250;
  wire [31:0] alu_0_i_y_out;
  wire alu_0_i_y2_out;
  wire [11:0] alu_0_i_y3_out;
  wire [31:0] n17257_o;
  wire [11:0] n17258_o;
  wire [11:0] n17259_o;
  wire [31:0] alu_1_i_n17260;
  wire alu_1_i_n17261;
  wire [11:0] alu_1_i_n17262;
  wire [31:0] alu_1_i_y_out;
  wire alu_1_i_y2_out;
  wire [11:0] alu_1_i_y3_out;
  wire [31:0] n17269_o;
  wire [11:0] n17270_o;
  wire [11:0] n17271_o;
  wire [31:0] alu_2_i_n17272;
  wire alu_2_i_n17273;
  wire [11:0] alu_2_i_n17274;
  wire [31:0] alu_2_i_y_out;
  wire alu_2_i_y2_out;
  wire [11:0] alu_2_i_y3_out;
  wire [31:0] n17281_o;
  wire [11:0] n17282_o;
  wire [11:0] n17283_o;
  wire [31:0] alu_3_i_n17284;
  wire alu_3_i_n17285;
  wire [11:0] alu_3_i_n17286;
  wire [31:0] alu_3_i_y_out;
  wire alu_3_i_y2_out;
  wire [11:0] alu_3_i_y3_out;
  wire [31:0] n17293_o;
  wire [11:0] n17294_o;
  wire [11:0] n17295_o;
  wire [31:0] alu_4_i_n17296;
  wire alu_4_i_n17297;
  wire [11:0] alu_4_i_n17298;
  wire [31:0] alu_4_i_y_out;
  wire alu_4_i_y2_out;
  wire [11:0] alu_4_i_y3_out;
  wire [31:0] n17305_o;
  wire [11:0] n17306_o;
  wire [11:0] n17307_o;
  wire [31:0] alu_5_i_n17308;
  wire alu_5_i_n17309;
  wire [11:0] alu_5_i_n17310;
  wire [31:0] alu_5_i_y_out;
  wire alu_5_i_y2_out;
  wire [11:0] alu_5_i_y3_out;
  wire [31:0] n17317_o;
  wire [11:0] n17318_o;
  wire [11:0] n17319_o;
  wire [31:0] alu_6_i_n17320;
  wire alu_6_i_n17321;
  wire [11:0] alu_6_i_n17322;
  wire [31:0] alu_6_i_y_out;
  wire alu_6_i_y2_out;
  wire [11:0] alu_6_i_y3_out;
  wire [31:0] n17329_o;
  wire [11:0] n17330_o;
  wire [11:0] n17331_o;
  wire [31:0] alu_7_i_n17332;
  wire alu_7_i_n17333;
  wire [11:0] alu_7_i_n17334;
  wire [31:0] alu_7_i_y_out;
  wire alu_7_i_y2_out;
  wire [11:0] alu_7_i_y3_out;
  wire n17341_o;
  wire n17342_o;
  wire [12:0] ialu_i_n17343;
  wire ialu_i_n17344;
  wire ialu_i_n17345;
  wire [12:0] ialu_i_y_out;
  wire ialu_i_y_neg_out;
  wire ialu_i_y_zero_out;
  wire [95:0] register_bank_i_n17354;
  wire [95:0] register_bank_i_n17355;
  wire [16:0] n17356_o;
  wire [16:0] n17357_o;
  wire [95:0] register_bank_i_n17358;
  wire register_bank_i_n17359;
  wire register_bank_i_n17360;
  wire [2:0] register_bank_i_n17361;
  wire [2:0] register_bank_i_n17362;
  wire [1:0] register_bank_i_n17363;
  wire [2:0] register_bank_i_n17364;
  wire [2:0] register_bank_i_n17365;
  wire register_bank_i_n17366;
  wire [1:0] register_bank_i_n17367;
  wire [1:0] register_bank_i_n17368;
  wire register_bank_i_n17369;
  wire [1:0] register_bank_i_n17370;
  wire register_bank_i_rd_en_out;
  wire [95:0] register_bank_i_rd_x1_data_out;
  wire [95:0] register_bank_i_rd_x2_data_out;
  wire [95:0] register_bank_i_dp_readdata_out;
  wire register_bank_i_dp_readdata_vm_out;
  wire register_bank_i_dp_readena_out;
  wire [2:0] register_bank_i_dp_read_vector_out;
  wire [2:0] register_bank_i_dp_read_vaddr_out;
  wire [1:0] register_bank_i_dp_read_scatter_out;
  wire [2:0] register_bank_i_dp_read_scatter_cnt_out;
  wire [2:0] register_bank_i_dp_read_scatter_vector_out;
  wire register_bank_i_dp_read_gen_valid_out;
  wire [1:0] register_bank_i_dp_read_data_flow_out;
  wire [1:0] register_bank_i_dp_read_data_type_out;
  wire register_bank_i_dp_read_stream_out;
  wire [1:0] register_bank_i_dp_read_stream_id_out;
  wire [4:0] instr_decoder2_i_n17403;
  wire instr_decoder2_i_n17404;
  wire [3:0] instr_decoder2_i_n17405;
  wire instr_decoder2_i_n17406;
  wire instr_decoder2_i_n17407;
  wire instr_decoder2_i_n17408;
  wire instr_decoder2_i_n17409;
  wire [11:0] instr_decoder2_i_n17410;
  wire [11:0] instr_decoder2_i_n17411;
  wire [11:0] instr_decoder2_i_n17412;
  wire instr_decoder2_i_n17413;
  wire instr_decoder2_i_n17414;
  wire instr_decoder2_i_n17415;
  wire [7:0] instr_decoder2_i_n17416;
  wire instr_decoder2_i_n17417;
  wire [11:0] instr_decoder2_i_n17418;
  wire instr_decoder2_i_n17419;
  wire instr_decoder2_i_n17420;
  wire [3:0] instr_decoder2_i_n17421;
  wire [3:0] instr_decoder2_i_n17422;
  wire instr_decoder2_i_n17423;
  wire instr_decoder2_i_n17424;
  wire [2:0] instr_decoder2_i_n17425;
  wire [12:0] instr_decoder2_i_n17426;
  wire instr_decoder2_i_n17427;
  wire [4:0] instr_decoder2_i_n17428;
  wire [12:0] instr_decoder2_i_n17429;
  wire [12:0] instr_decoder2_i_n17430;
  wire [7:0] instr_decoder2_i_n17431;
  wire [7:0] instr_decoder2_i_n17432;
  wire [4:0] instr_decoder2_i_opcode1_out;
  wire instr_decoder2_i_en1_out;
  wire [3:0] instr_decoder2_i_instruction_tid_out;
  wire instr_decoder2_i_xreg1_out;
  wire instr_decoder2_i_flag1_out;
  wire instr_decoder2_i_wren_out;
  wire instr_decoder2_i_vm_out;
  wire [11:0] instr_decoder2_i_x1_addr1_out;
  wire [11:0] instr_decoder2_i_x2_addr1_out;
  wire [11:0] instr_decoder2_i_y_addr1_out;
  wire instr_decoder2_i_x1_vector_out;
  wire instr_decoder2_i_x2_vector_out;
  wire instr_decoder2_i_y_vector_out;
  wire [7:0] instr_decoder2_i_vector_lane_out;
  wire instr_decoder2_i_x1_c1_en_out;
  wire [11:0] instr_decoder2_i_x1_c1_out;
  wire instr_decoder2_i_i_rd_en_out;
  wire instr_decoder2_i_i_rd_vm_out;
  wire [3:0] instr_decoder2_i_i_rd_tid_out;
  wire [3:0] instr_decoder2_i_i_wr_tid_out;
  wire instr_decoder2_i_i_wr_en_out;
  wire instr_decoder2_i_i_wr_vm_out;
  wire [2:0] instr_decoder2_i_i_wr_addr_out;
  wire [12:0] instr_decoder2_i_i_wr_data_out;
  wire instr_decoder2_i_wr_lane_out;
  wire [4:0] instr_decoder2_i_i_opcode_out;
  wire [12:0] instr_decoder2_i_i_x1_out;
  wire [12:0] instr_decoder2_i_i_x2_out;
  wire [7:0] instr_decoder2_i_result_waddr_out;
  wire [7:0] instr_decoder2_i_result_raddr_out;
  wire instr_dispatch2_i1_n17493;
  wire instr_dispatch2_i1_n17494;
  wire [11:0] instr_dispatch2_i1_n17495;
  wire [11:0] instr_dispatch2_i1_n17496;
  wire instr_dispatch2_i1_n17497;
  wire instr_dispatch2_i1_n17498;
  wire instr_dispatch2_i1_n17499;
  wire instr_dispatch2_i1_n17500;
  wire instr_dispatch2_i1_n17501;
  wire instr_dispatch2_i1_n17502;
  wire instr_dispatch2_i1_n17503;
  wire instr_dispatch2_i1_n17504;
  wire [11:0] instr_dispatch2_i1_n17505;
  wire [7:0] instr_dispatch2_i1_n17506;
  wire [95:0] instr_dispatch2_i1_n17507;
  wire [7:0] instr_dispatch2_i1_n17508;
  wire [95:0] instr_dispatch2_i1_n17509;
  wire [95:0] instr_dispatch2_i1_n17510;
  wire [11:0] instr_dispatch2_i1_n17511;
  wire [4:0] instr_dispatch2_i1_n17512;
  wire [3:0] instr_dispatch2_i1_n17513;
  wire instr_dispatch2_i1_rd_en_out;
  wire instr_dispatch2_i1_rd_vm_out;
  wire [11:0] instr_dispatch2_i1_rd_x1_addr_out;
  wire [11:0] instr_dispatch2_i1_rd_x2_addr_out;
  wire instr_dispatch2_i1_rd_x1_vector_out;
  wire instr_dispatch2_i1_rd_x2_vector_out;
  wire instr_dispatch2_i1_wr_xreg_out;
  wire instr_dispatch2_i1_wr_flag_out;
  wire instr_dispatch2_i1_wr_xreg_flag_out;
  wire instr_dispatch2_i1_wr_en_out;
  wire instr_dispatch2_i1_wr_vm_out;
  wire instr_dispatch2_i1_wr_vector_out;
  wire [11:0] instr_dispatch2_i1_wr_addr_out;
  wire [7:0] instr_dispatch2_i1_wr_result_addr_out;
  wire [95:0] instr_dispatch2_i1_wr_data_out;
  wire [7:0] instr_dispatch2_i1_wr_lane_out;
  wire [95:0] instr_dispatch2_i1_mu_x1_out;
  wire [95:0] instr_dispatch2_i1_mu_x2_out;
  wire [11:0] instr_dispatch2_i1_mu_x_scalar_out;
  wire [4:0] instr_dispatch2_i1_mu_opcode_out;
  wire [3:0] instr_dispatch2_i1_mu_tid_out;
  wire [255:0] n17559_o;
  wire [95:0] n17560_o;
  wire [7:0] n17561_o;
  wire [95:0] n17562_o;
  reg [95:0] n17563_q;
  wire [95:0] n17564_o;
  reg [95:0] n17565_q;
  reg n17566_q;
  reg n17567_q;
  wire n17568_o;
  reg n17569_q;
  wire [1:0] n17570_o;
  reg [1:0] n17571_q;
  wire [1:0] n17572_o;
  reg [1:0] n17573_q;
  wire [2:0] n17574_o;
  reg [2:0] n17575_q;
  wire [2:0] n17576_o;
  reg [2:0] n17577_q;
  wire n17578_o;
  reg n17579_q;
  wire [1:0] n17580_o;
  reg [1:0] n17581_q;
  reg [2:0] n17582_q;
  reg [2:0] n17583_q;
  reg [1:0] n17584_q;
  reg [2:0] n17587_q;
  reg [2:0] n17588_q;
  reg n17589_q;
  reg [1:0] n17590_q;
  reg [1:0] n17591_q;
  reg n17592_q;
  reg [1:0] n17593_q;
  reg [21:0] n17594_q;
  reg [2:0] n17595_q;
  reg [21:0] n17596_q;
  reg [95:0] n17597_q;
  wire n17598_o;
  reg n17599_q;
  wire n17600_o;
  reg n17601_q;
  wire n17602_o;
  reg n17603_q;
  reg [21:0] n17606_q;
  reg [21:0] n17607_q;
  wire [5:0] n17608_o;
  reg [5:0] n17609_q;
  wire n17610_o;
  reg n17611_q;
  wire [2:0] n17614_o;
  reg [2:0] n17615_q;
  wire [1:0] n17616_o;
  reg [1:0] n17617_q;
  wire n17618_o;
  reg n17619_q;
  wire [21:0] n17620_o;
  reg [21:0] n17621_q;
  wire n17622_o;
  reg n17623_q;
  wire [2:0] n17624_o;
  reg [2:0] n17625_q;
  wire [1:0] n17626_o;
  reg [1:0] n17627_q;
  wire n17628_o;
  wire n17629_o;
  wire n17630_o;
  reg n17631_q;
  wire n17632_o;
  wire n17633_o;
  wire [21:0] n17634_o;
  reg [21:0] n17635_q;
  wire n17636_o;
  reg n17637_q;
  wire [1:0] n17638_o;
  reg [1:0] n17639_q;
  wire [1:0] n17640_o;
  reg [1:0] n17641_q;
  wire n17642_o;
  reg n17643_q;
  wire [1:0] n17644_o;
  reg [1:0] n17645_q;
  reg [83:0] n17646_q;
  wire [95:0] n17647_o;
  reg [2:0] n17648_q;
  reg [2:0] n17649_q;
  reg [2:0] n17650_q;
  reg [79:0] n17652_q;
  reg [31:0] n17653_q;
  reg n17654_q;
  reg n17655_q;
  reg n17656_q;
  reg [1:0] n17657_q;
  reg [3:0] n17658_q;
  reg n17659_q;
  reg [3:0] n17660_q;
  reg n17661_q;
  reg [3:0] n17662_q;
  reg n17663_q;
  reg n17664_q;
  reg [1:0] n17665_q;
  reg [27:0] n17666_q;
  reg n17667_q;
  reg n17668_q;
  reg n17670_q;
  reg n17671_q;
  reg n17673_q;
  reg n17674_q;
  reg n17675_q;
  reg [21:0] n17676_q;
  reg n17677_q;
  reg [21:0] n17678_q;
  reg [21:0] n17679_q;
  reg n17680_q;
  reg [21:0] n17681_q;
  reg [5:0] n17682_q;
  reg n17683_q;
  reg n17684_q;
  reg n17685_q;
  reg [2:0] n17686_q;
  reg [1:0] n17687_q;
  reg n17688_q;
  reg n17689_q;
  reg [2:0] n17690_q;
  reg [1:0] n17691_q;
  reg n17692_q;
  reg [1:0] n17693_q;
  reg [1:0] n17694_q;
  reg n17695_q;
  reg [1:0] n17696_q;
  reg [95:0] n17697_q;
  reg n17698_q;
  wire [2:0] n17699_o;
  wire [2:0] n17700_o;
  assign i_y_neg_out = n17341_o;
  assign i_y_zero_out = n17342_o;
  assign dp_readdata_out = n17014_o;
  assign dp_readdata_vm_out = n17016_o;
  assign dp_readena_out = dp_readena_r;
  assign dp_read_vector_out = n17699_o;
  assign dp_read_vaddr_out = n17700_o;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_r;
  assign dp_read_data_flow_out = n16994_o;
  assign dp_read_data_type_out = n16996_o;
  assign dp_read_stream_out = n16998_o;
  assign dp_read_stream_id_out = n17000_o;
  /* ../../HW/src/pcore/pcore.vhd:88:8  */
  assign rd_x1_data1 = register_bank_i_n17354; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:89:8  */
  assign rd_x2_data1 = register_bank_i_n17355; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:90:8  */
  assign rd_en1 = instr_dispatch2_i1_n17493; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:91:8  */
  assign rd_vm = instr_dispatch2_i1_n17494; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:92:8  */
  assign wr_en1 = instr_dispatch2_i1_n17502; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:93:8  */
  assign wr_xreg1 = instr_dispatch2_i1_n17499; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:94:8  */
  assign wr_flag1 = instr_dispatch2_i1_n17500; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:95:8  */
  assign wr_xreg_flag1 = instr_dispatch2_i1_n17501; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:96:8  */
  assign wr_data1 = instr_dispatch2_i1_n17507; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:97:8  */
  assign wr_vector_lane = instr_dispatch2_i1_n17508; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:98:8  */
  assign x1_addr1 = instr_decoder2_i_n17410; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:99:8  */
  assign x2_addr1 = instr_decoder2_i_n17411; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:100:8  */
  assign y_addr1 = instr_decoder2_i_n17412; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:101:8  */
  assign rd_lane = iregister_i_n17192; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:102:8  */
  assign wr_lane = instr_decoder2_i_n17427; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:103:8  */
  assign opcode1 = instr_decoder2_i_n17403; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:107:8  */
  assign mu_x1 = instr_dispatch2_i1_n17509; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:108:8  */
  assign mu_x2 = instr_dispatch2_i1_n17510; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:109:8  */
  assign mu_x_scalar = instr_dispatch2_i1_n17511; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:110:8  */
  assign mu_y = n17559_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:111:8  */
  assign mu_y2 = n17560_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:112:8  */
  assign mu_result = n17561_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:113:8  */
  assign mu_opcodes = instr_dispatch2_i1_n17512; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:114:8  */
  assign mu_tid = instr_dispatch2_i1_n17513; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:115:8  */
  assign tid_decoder2dispatch = instr_decoder2_i_n17405; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:117:8  */
  assign write = n17242_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:118:8  */
  assign read = n17215_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:120:8  */
  assign dp_mcast_addr = n17008_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:122:8  */
  assign rd_x1_addr1 = instr_dispatch2_i1_n17495; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:123:8  */
  assign rd_x2_addr1 = instr_dispatch2_i1_n17496; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:124:8  */
  assign wr_addr1 = instr_dispatch2_i1_n17505; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:125:8  */
  assign wr_result_addr1 = instr_dispatch2_i1_n17506; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:127:8  */
  assign dp_rd_pid = n17006_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:128:8  */
  assign dp_rd_cid = n17007_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:129:8  */
  assign en1 = instr_decoder2_i_n17404; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:130:8  */
  assign mu_vm = instr_decoder2_i_n17409; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:131:8  */
  assign mu_xreg1 = instr_decoder2_i_n17406; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:132:8  */
  assign mu_flag1 = instr_decoder2_i_n17407; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:133:8  */
  assign mu_wren = instr_decoder2_i_n17408; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:136:8  */
  assign x1_c1_en = instr_decoder2_i_n17417; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:137:8  */
  assign x1_c1 = instr_decoder2_i_n17418; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:140:8  */
  assign x1_vector = instr_decoder2_i_n17413; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:141:8  */
  assign x2_vector = instr_decoder2_i_n17414; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:142:8  */
  assign y_vector = instr_decoder2_i_n17415; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:143:8  */
  assign vector_lane = instr_decoder2_i_n17416; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:144:8  */
  assign rd_x1_vector1 = instr_dispatch2_i1_n17497; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:145:8  */
  assign rd_x2_vector1 = instr_dispatch2_i1_n17498; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:146:8  */
  assign wr_vector = instr_dispatch2_i1_n17504; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:149:8  */
  assign i_rd_en1 = instr_decoder2_i_n17419; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:150:8  */
  assign i_rd_vm = instr_decoder2_i_n17420; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:151:8  */
  assign i_rd_tid1 = instr_decoder2_i_n17421; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:152:8  */
  assign i_rd_data1 = iregister_i_n17191; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:153:8  */
  assign i_wr_tid1 = instr_decoder2_i_n17422; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:154:8  */
  assign i_wr_en1 = instr_decoder2_i_n17423; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:155:8  */
  assign i_wr_vm = instr_decoder2_i_n17424; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:156:8  */
  assign i_wr_addr1 = instr_decoder2_i_n17425; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:157:8  */
  assign i_wr_data1 = instr_decoder2_i_n17426; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:159:8  */
  assign dp_readdata_r = n17563_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:160:8  */
  assign dp_readdata2_r = n17565_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:161:8  */
  assign dp_readena_r = n17566_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:162:8  */
  assign dp_readdata_vm_r = n17567_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:163:8  */
  assign dp_read_gen_valid2_r = n17569_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:164:8  */
  assign dp_read_data_flow2_r = n17571_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:165:8  */
  assign dp_read_data_type2_r = n17573_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:166:8  */
  assign dp_read_vector2_r = n17575_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:167:8  */
  assign dp_read_vaddr2_r = n17577_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:168:8  */
  assign dp_read_stream2_r = n17579_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:169:8  */
  assign dp_read_stream_id2_r = n17581_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:173:8  */
  assign i_opcode = instr_decoder2_i_n17428; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:174:8  */
  assign i_x1 = instr_decoder2_i_n17429; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:175:8  */
  assign i_x2 = instr_decoder2_i_n17430; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:176:8  */
  assign i_y = ialu_i_n17343; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:177:8  */
  assign i_y_neg = ialu_i_n17344; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:178:8  */
  assign i_y_zero = ialu_i_n17345; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:180:8  */
  assign wr_vm = instr_dispatch2_i1_n17503; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:181:8  */
  assign result_write_addr = wr_result_addr1; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:183:8  */
  assign result_raddr1 = instr_decoder2_i_n17431; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:184:8  */
  assign result_waddr1 = instr_decoder2_i_n17432; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:185:8  */
  assign result_read = xregister_file_i_n17185; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:186:8  */
  assign xreg_read = xregister_file_i_n17186; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:188:8  */
  assign dp_rd_vm = n16674_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:189:8  */
  assign dp_rd_fork = n16675_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:190:8  */
  assign dp_wr_vm = n16714_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:192:8  */
  assign dp_rd_addr = n16676_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:193:8  */
  assign dp_wr_addr = n16716_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:194:8  */
  assign dp_wr_mcast = n16717_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:195:8  */
  assign dp_write = n16718_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:196:8  */
  assign dp_write_vector = n16719_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:197:8  */
  assign dp_write_scatter = n16720_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:198:8  */
  assign dp_write_share = n16721_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:199:8  */
  assign dp_write_step = n16722_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:201:8  */
  assign dp_read = n16677_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:202:8  */
  assign dp_read_vector = n16678_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:203:8  */
  assign dp_read_scatter = n16679_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:204:8  */
  assign dp_read_share = n16680_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:205:8  */
  assign dp_read_step = n16681_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:206:8  */
  assign dp_read_gen_valid = n16682_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:207:8  */
  assign dp_read_data_flow = n16683_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:208:8  */
  assign dp_read_data_type = n16684_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:209:8  */
  assign dp_read_stream = n16685_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:210:8  */
  assign dp_read_stream_id = n16686_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:211:8  */
  assign dp_writedata = n16968_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_cnt = n16687_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:600:10  */
  assign read_scatter_vector = n16688_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:214:8  */
  assign write_scatter_cnt = n16724_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:216:8  */
  assign write_scatter_curr = n16727_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:217:8  */
  assign write_scatter_curr_r = n17582_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:219:8  */
  assign gen_read_vector_r = n17583_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:220:8  */
  assign gen_read_scatter_r = n17584_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:223:8  */
  assign gen_read_scatter_cnt_r = n17587_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:224:8  */
  assign gen_read_scatter_vector_r = n17588_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:225:8  */
  assign gen_read_gen_valid_r = n17589_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:226:8  */
  assign gen_read_data_flow_r = n17590_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:227:8  */
  assign gen_read_data_type_r = n17591_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:228:8  */
  assign gen_read_stream_r = n17592_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:229:8  */
  assign gen_read_stream_id_r = n17593_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:230:8  */
  assign gen_rd_addr_r = n17594_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:231:8  */
  assign gen_write_vector_r = n17595_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:232:8  */
  assign gen_wr_addr_r = n17596_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:233:8  */
  assign gen_writedata_r = n17597_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:235:8  */
  assign dp_rd_vm_r = n17599_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:236:8  */
  assign dp_rd_fork_r = n17601_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:237:8  */
  assign dp_wr_vm_r = n17603_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:239:8  */
  assign dp_rd_addr_r = n17606_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:240:8  */
  assign dp_wr_addr_r = n17607_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:241:8  */
  assign dp_wr_mcast_r = n17609_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:242:8  */
  assign dp_write_r = n17611_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:244:8  */
  assign dp_write_vector_r = n17615_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:245:8  */
  assign dp_write_scatter_r = n17617_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:246:8  */
  assign dp_write_share_r = n17619_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:247:8  */
  assign dp_write_step_r = n17621_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:248:8  */
  assign dp_read_r = n17623_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:249:8  */
  assign dp_read_vector_r = n17625_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:250:8  */
  assign dp_read_scatter_r = n17627_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:251:8  */
  assign dp_read_share_r = n17631_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:252:8  */
  assign dp_read_step_r = n17635_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:253:8  */
  assign dp_read_gen_valid_r = n17637_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:254:8  */
  assign dp_read_data_flow_r = n17639_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:255:8  */
  assign dp_read_data_type_r = n17641_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:256:8  */
  assign dp_read_stream_r = n17643_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:257:8  */
  assign dp_read_stream_id_r = n17645_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:258:8  */
  assign dp_writedata_r = n17647_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:259:8  */
  assign read_scatter_cnt_r = n17648_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:260:8  */
  assign read_scatter_vector_r = n17649_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:261:8  */
  assign write_scatter_cnt_r = n17650_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:264:8  */
  assign read_match = n16992_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:265:8  */
  assign write_match = n16653_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:267:8  */
  assign dp_readena_vm = register_bank_i_n17360; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:269:8  */
  assign dp_read_vector_vm = register_bank_i_n17361; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:271:8  */
  assign dp_read_vaddr_vm = register_bank_i_n17362; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:273:8  */
  assign dp_read_scatter_vm = register_bank_i_n17363; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:274:8  */
  assign dp_read_scatter_cnt_vm = register_bank_i_n17364; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:275:8  */
  assign dp_read_scatter_vector_vm = register_bank_i_n17365; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:276:8  */
  assign dp_readdata_vm = register_bank_i_n17358; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:277:8  */
  assign dp_readdata_vm_vm = register_bank_i_n17359; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:278:8  */
  assign dp_read_gen_valid_vm = register_bank_i_n17366; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:279:8  */
  assign dp_read_data_flow_vm = register_bank_i_n17367; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:280:8  */
  assign dp_read_data_type_vm = register_bank_i_n17368; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:281:8  */
  assign dp_read_stream_vm = register_bank_i_n17369; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:282:8  */
  assign dp_read_stream_id_vm = register_bank_i_n17370; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:284:8  */
  assign tid_valid1 = n16531_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:285:8  */
  assign pre_tid_valid1 = n16532_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:286:8  */
  assign pre_pre_tid_valid1 = n16533_o; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:288:8  */
  assign instruction_mu_r = n17652_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:289:8  */
  assign instruction_imu_r = n17653_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:290:8  */
  assign instruction_mu_valid_r = n17654_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:291:8  */
  assign instruction_imu_valid_r = n17655_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:293:8  */
  assign vm_r = n17656_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:294:8  */
  assign data_model_r = n17657_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:295:8  */
  assign tid_r = n17658_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:296:8  */
  assign tid_valid1_r = n17659_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:297:8  */
  assign pre_tid_r = n17660_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:298:8  */
  assign pre_tid_valid1_r = n17661_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:299:8  */
  assign pre_pre_tid_r = n17662_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:300:8  */
  assign pre_pre_tid_valid1_r = n17663_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:301:8  */
  assign pre_pre_vm_r = n17664_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:302:8  */
  assign pre_pre_data_model_r = n17665_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:303:8  */
  assign pre_iregister_auto_r = n17666_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:305:8  */
  assign gen_write_r = n17667_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:306:8  */
  assign gen_write_vm_r = n17668_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:308:8  */
  assign gen_read_r = n17670_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:309:8  */
  assign gen_read_vm_r = n17671_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:312:8  */
  assign dp_rd_vm_in_r = n17673_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:313:8  */
  assign dp_wr_vm_in_r = n17674_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:314:8  */
  assign dp_code_in_r = n17675_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:315:8  */
  assign dp_rd_addr_in_r = n17676_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:316:8  */
  assign dp_rd_share_in_r = n17677_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:317:8  */
  assign dp_rd_step_in_r = n17678_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:318:8  */
  assign dp_wr_addr_in_r = n17679_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:319:8  */
  assign dp_wr_share_in_r = n17680_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:320:8  */
  assign dp_wr_step_in_r = n17681_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:321:8  */
  assign dp_wr_mcast_in_r = n17682_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:322:8  */
  assign dp_write_in_r = n17683_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:323:8  */
  assign dp_wr_fork_in_r = n17684_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:324:8  */
  assign dp_write_gen_valid_in_r = n17685_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:325:8  */
  assign dp_write_vector_in_r = n17686_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:326:8  */
  assign dp_write_scatter_in_r = n17687_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:327:8  */
  assign dp_rd_fork_in_r = n17688_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:328:8  */
  assign dp_read_in_r = n17689_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:329:8  */
  assign dp_read_vector_in_r = n17690_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:330:8  */
  assign dp_read_scatter_in_r = n17691_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:331:8  */
  assign dp_read_gen_valid_in_r = n17692_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:332:8  */
  assign dp_read_data_flow_in_r = n17693_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:333:8  */
  assign dp_read_data_type_in_r = n17694_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:334:8  */
  assign dp_read_stream_in_r = n17695_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:335:8  */
  assign dp_read_stream_id_in_r = n17696_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:336:8  */
  assign dp_writedata_in_r = n17697_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:337:8  */
  assign dp_config_in_r = n17698_q; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:341:28  */
  assign n16531_o = tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:343:36  */
  assign n16532_o = pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:345:44  */
  assign n16533_o = pre_pre_tid_valid1_r & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:349:13  */
  assign n16536_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:423:31  */
  assign n16624_o = dp_wr_mcast_in_r[4:0];
  /* ../../HW/src/pcore/pcore.vhd:424:36  */
  assign n16625_o = dp_wr_mcast_in_r[5];
  /* ../../HW/src/pcore/pcore.vhd:425:35  */
  assign n16626_o = dp_wr_addr_in_r[16:12];
  /* ../../HW/src/pcore/pcore.vhd:426:22  */
  assign n16627_o = ~dp_wr_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:426:4  */
  assign n16630_o = n16627_o ? 3'b000 : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:432:56  */
  assign n16632_o = n16626_o + n16624_o;
  /* ../../HW/src/pcore/pcore.vhd:433:44  */
  assign n16633_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:27  */
  assign n16634_o = n16633_o & dp_write_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:69  */
  assign n16635_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:433:50  */
  assign n16636_o = n16635_o & n16634_o;
  /* ../../HW/src/pcore/pcore.vhd:435:38  */
  assign n16637_o = n16624_o & n16626_o;
  assign n16638_o = {n16630_o, 2'b00};
  /* ../../HW/src/pcore/pcore.vhd:435:65  */
  assign n16639_o = n16624_o & n16638_o;
  /* ../../HW/src/pcore/pcore.vhd:435:55  */
  assign n16640_o = n16637_o == n16639_o;
  /* ../../HW/src/pcore/pcore.vhd:435:25  */
  assign n16641_o = n16640_o & n16625_o;
  /* ../../HW/src/pcore/pcore.vhd:437:20  */
  assign n16642_o = ~n16625_o;
  assign n16643_o = {n16630_o, 2'b00};
  /* ../../HW/src/pcore/pcore.vhd:437:49  */
  assign n16644_o = $unsigned(n16643_o) >= $unsigned(n16626_o);
  /* ../../HW/src/pcore/pcore.vhd:437:25  */
  assign n16645_o = n16644_o & n16642_o;
  assign n16646_o = {n16630_o, 2'b00};
  /* ../../HW/src/pcore/pcore.vhd:437:100  */
  assign n16647_o = $unsigned(n16646_o) <= $unsigned(n16632_o);
  /* ../../HW/src/pcore/pcore.vhd:437:76  */
  assign n16648_o = n16647_o & n16645_o;
  /* ../../HW/src/pcore/pcore.vhd:436:7  */
  assign n16649_o = n16641_o | n16648_o;
  /* ../../HW/src/pcore/pcore.vhd:433:75  */
  assign n16650_o = n16649_o & n16636_o;
  /* ../../HW/src/pcore/pcore.vhd:433:4  */
  assign n16653_o = n16650_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:461:24  */
  assign n16659_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:467:27  */
  assign n16661_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:467:4  */
  assign n16663_o = n16661_o ? 3'b000 : dp_read_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:481:47  */
  assign n16665_o = dp_read_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:481:23  */
  assign n16666_o = n16665_o & read_match;
  /* ../../HW/src/pcore/pcore.vhd:481:64  */
  assign n16667_o = dp_read_gen_valid_in_r & n16666_o;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n16669_o = n16667_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:481:4  */
  assign n16671_o = n16667_o ? dp_read_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:504:42  */
  assign n16673_o = read_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16674_o = n16659_o ? dp_rd_vm_in_r : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16675_o = n16659_o ? dp_rd_fork_in_r : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16676_o = n16659_o ? dp_rd_addr_in_r : dp_rd_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16677_o = n16659_o ? dp_read_in_r : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16678_o = n16659_o ? n16663_o : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16679_o = n16659_o ? dp_read_scatter_in_r : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16680_o = n16659_o ? dp_rd_share_in_r : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16681_o = n16659_o ? dp_rd_step_in_r : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16682_o = n16659_o ? dp_read_gen_valid_in_r : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16683_o = n16659_o ? dp_read_data_flow_in_r : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16684_o = n16659_o ? dp_read_data_type_in_r : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16685_o = n16659_o ? dp_read_stream_in_r : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16686_o = n16659_o ? dp_read_stream_id_in_r : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16687_o = n16659_o ? n16669_o : n16673_o;
  /* ../../HW/src/pcore/pcore.vhd:461:1  */
  assign n16688_o = n16659_o ? n16671_o : read_scatter_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:24  */
  assign n16693_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:526:35  */
  assign n16694_o = ~dp_code_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:30  */
  assign n16695_o = dp_write_in_r & n16694_o;
  /* ../../HW/src/pcore/pcore.vhd:526:58  */
  assign n16696_o = ~dp_config_in_r;
  /* ../../HW/src/pcore/pcore.vhd:526:53  */
  assign n16697_o = n16695_o & n16696_o;
  /* ../../HW/src/pcore/pcore.vhd:527:28  */
  assign n16699_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:527:4  */
  assign n16701_o = n16699_o ? 3'b000 : dp_write_vector_in_r;
  /* ../../HW/src/pcore/pcore.vhd:536:49  */
  assign n16703_o = dp_write_scatter_in_r != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:536:24  */
  assign n16704_o = n16703_o & write_match;
  /* ../../HW/src/pcore/pcore.vhd:536:66  */
  assign n16705_o = dp_write_gen_valid_in_r & n16704_o;
  /* ../../HW/src/pcore/pcore.vhd:536:4  */
  assign n16707_o = n16705_o ? dp_write_vector_in_r : 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:557:44  */
  assign n16711_o = write_scatter_cnt_r - 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:559:46  */
  assign n16713_o = write_scatter_curr_r + 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16714_o = n16693_o ? dp_wr_vm_in_r : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16716_o = n16693_o ? dp_wr_addr_in_r : dp_wr_addr_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16717_o = n16693_o ? dp_wr_mcast_in_r : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16718_o = n16693_o ? n16697_o : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16719_o = n16693_o ? n16701_o : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16720_o = n16693_o ? dp_write_scatter_in_r : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16721_o = n16693_o ? dp_wr_share_in_r : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16722_o = n16693_o ? dp_wr_step_in_r : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16724_o = n16693_o ? n16707_o : n16711_o;
  /* ../../HW/src/pcore/pcore.vhd:520:1  */
  assign n16727_o = n16693_o ? 3'b000 : n16713_o;
  /* ../../HW/src/pcore/pcore.vhd:573:16  */
  assign n16732_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:590:28  */
  assign n16735_o = dp_read_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:591:29  */
  assign n16736_o = ~dp_read_share;
  /* ../../HW/src/pcore/pcore.vhd:592:46  */
  assign n16737_o = dp_rd_addr + dp_read_step;
  /* ../../HW/src/pcore/pcore.vhd:594:46  */
  assign n16739_o = dp_rd_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:591:13  */
  assign n16740_o = n16736_o ? n16737_o : n16739_o;
  /* ../../HW/src/pcore/pcore.vhd:597:43  */
  assign n16742_o = dp_rd_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:590:10  */
  assign n16743_o = n16735_o ? n16740_o : n16742_o;
  /* ../../HW/src/pcore/pcore.vhd:600:32  */
  assign n16745_o = read_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:630:16  */
  assign n16809_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:690:16  */
  assign n16878_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:707:29  */
  assign n16881_o = dp_write_scatter == 2'b01;
  /* ../../HW/src/pcore/pcore.vhd:708:30  */
  assign n16882_o = ~dp_write_share;
  /* ../../HW/src/pcore/pcore.vhd:709:46  */
  assign n16883_o = dp_wr_addr + dp_write_step;
  /* ../../HW/src/pcore/pcore.vhd:711:46  */
  assign n16885_o = dp_wr_addr - 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:708:13  */
  assign n16886_o = n16882_o ? n16883_o : n16885_o;
  /* ../../HW/src/pcore/pcore.vhd:714:43  */
  assign n16888_o = dp_wr_addr + 22'b0000000000000000001000;
  /* ../../HW/src/pcore/pcore.vhd:707:10  */
  assign n16889_o = n16881_o ? n16886_o : n16888_o;
  /* ../../HW/src/pcore/pcore.vhd:717:33  */
  assign n16891_o = write_scatter_cnt_r == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:728:96  */
  assign n16892_o = dp_writedata_in_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:731:93  */
  assign n16893_o = dp_writedata_r[95:12];
  /* ../../HW/src/pcore/pcore.vhd:717:10  */
  assign n16903_o = n16891_o ? n16892_o : n16893_o;
  assign n16945_o = dp_writedata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n16946_o = n16878_o ? 12'b000000000000 : n16945_o;
  /* ../../HW/src/pcore/pcore.vhd:748:20  */
  assign n16960_o = dp_write_scatter != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:750:12  */
  assign n16962_o = write_scatter_curr == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:751:69  */
  assign n16963_o = dp_writedata_in_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:753:66  */
  assign n16964_o = dp_writedata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:750:4  */
  assign n16965_o = n16962_o ? n16963_o : n16964_o;
  assign n16967_o = {84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000, n16965_o};
  /* ../../HW/src/pcore/pcore.vhd:748:1  */
  assign n16968_o = n16960_o ? n16967_o : dp_writedata_in_r;
  /* ../../HW/src/pcore/pcore.vhd:769:34  */
  assign n16974_o = dp_rd_addr_in_r[13:12];
  /* ../../HW/src/pcore/pcore.vhd:770:34  */
  assign n16975_o = dp_rd_addr_in_r[16:14];
  /* ../../HW/src/pcore/pcore.vhd:771:19  */
  assign n16976_o = ~dp_rd_fork_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:34  */
  assign n16978_o = n16974_o == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:772:25  */
  assign n16979_o = n16978_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:772:74  */
  assign n16981_o = n16975_o == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:772:65  */
  assign n16982_o = n16981_o & n16979_o;
  /* ../../HW/src/pcore/pcore.vhd:772:4  */
  assign n16985_o = n16982_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:778:34  */
  assign n16987_o = n16974_o == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:778:25  */
  assign n16988_o = n16987_o & dp_read_in_r;
  /* ../../HW/src/pcore/pcore.vhd:778:4  */
  assign n16991_o = n16988_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:771:1  */
  assign n16992_o = n16976_o ? n16985_o : n16991_o;
  /* ../../HW/src/pcore/pcore.vhd:792:47  */
  assign n16994_o = dp_readena_r ? dp_read_data_flow2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:793:47  */
  assign n16996_o = dp_readena_r ? dp_read_data_type2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:794:41  */
  assign n16998_o = dp_readena_r ? dp_read_stream2_r : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:795:47  */
  assign n17000_o = dp_readena_r ? dp_read_stream_id2_r : 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:798:33  */
  assign n17006_o = dp_rd_addr[13:12];
  /* ../../HW/src/pcore/pcore.vhd:799:33  */
  assign n17007_o = dp_rd_addr[16:14];
  /* ../../HW/src/pcore/pcore.vhd:800:28  */
  assign n17008_o = dp_wr_addr[16:12];
  /* ../../HW/src/pcore/pcore.vhd:808:16  */
  assign n17011_o = ~dp_readena_r;
  /* ../../HW/src/pcore/pcore.vhd:812:4  */
  assign n17012_o = dp_read_gen_valid2_r ? dp_readdata_r : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n17014_o = n17011_o ? 96'bZ : n17012_o;
  /* ../../HW/src/pcore/pcore.vhd:808:1  */
  assign n17016_o = n17011_o ? 1'bZ : dp_readdata_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:825:16  */
  assign n17021_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:870:16  */
  assign n17072_o = ~reset_in;
  /* ../../HW/src/pcore/pcore.vhd:886:38  */
  assign n17075_o = dp_read_scatter_vm != 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:887:54  */
  assign n17076_o = dp_read_scatter_vector_vm - dp_read_scatter_cnt_vm;
  /* ../../HW/src/pcore/pcore.vhd:891:105  */
  assign n17077_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:890:23  */
  assign n17079_o = n17076_o == 3'b111;
  /* ../../HW/src/pcore/pcore.vhd:893:105  */
  assign n17080_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:892:23  */
  assign n17082_o = n17076_o == 3'b110;
  /* ../../HW/src/pcore/pcore.vhd:895:105  */
  assign n17083_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:894:23  */
  assign n17085_o = n17076_o == 3'b101;
  /* ../../HW/src/pcore/pcore.vhd:897:105  */
  assign n17086_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:896:23  */
  assign n17088_o = n17076_o == 3'b100;
  /* ../../HW/src/pcore/pcore.vhd:899:105  */
  assign n17089_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:898:23  */
  assign n17091_o = n17076_o == 3'b011;
  /* ../../HW/src/pcore/pcore.vhd:901:105  */
  assign n17092_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:900:23  */
  assign n17094_o = n17076_o == 3'b010;
  /* ../../HW/src/pcore/pcore.vhd:903:105  */
  assign n17095_o = dp_readdata_vm[11:0];
  /* ../../HW/src/pcore/pcore.vhd:902:23  */
  assign n17097_o = n17076_o == 3'b001;
  /* ../../HW/src/pcore/pcore.vhd:905:105  */
  assign n17098_o = dp_readdata_vm[11:0];
  assign n17099_o = {n17097_o, n17094_o, n17091_o, n17088_o, n17085_o, n17082_o, n17079_o};
  assign n17100_o = dp_readdata_r[11:0];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17101_o = n17100_o;
      7'b0100000: n17101_o = n17100_o;
      7'b0010000: n17101_o = n17100_o;
      7'b0001000: n17101_o = n17100_o;
      7'b0000100: n17101_o = n17100_o;
      7'b0000010: n17101_o = n17100_o;
      7'b0000001: n17101_o = n17100_o;
      default: n17101_o = n17098_o;
    endcase
  assign n17102_o = dp_readdata_r[23:12];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17103_o = n17095_o;
      7'b0100000: n17103_o = n17102_o;
      7'b0010000: n17103_o = n17102_o;
      7'b0001000: n17103_o = n17102_o;
      7'b0000100: n17103_o = n17102_o;
      7'b0000010: n17103_o = n17102_o;
      7'b0000001: n17103_o = n17102_o;
      default: n17103_o = n17102_o;
    endcase
  assign n17104_o = dp_readdata_r[35:24];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17105_o = n17104_o;
      7'b0100000: n17105_o = n17092_o;
      7'b0010000: n17105_o = n17104_o;
      7'b0001000: n17105_o = n17104_o;
      7'b0000100: n17105_o = n17104_o;
      7'b0000010: n17105_o = n17104_o;
      7'b0000001: n17105_o = n17104_o;
      default: n17105_o = n17104_o;
    endcase
  assign n17106_o = dp_readdata_r[47:36];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17107_o = n17106_o;
      7'b0100000: n17107_o = n17106_o;
      7'b0010000: n17107_o = n17089_o;
      7'b0001000: n17107_o = n17106_o;
      7'b0000100: n17107_o = n17106_o;
      7'b0000010: n17107_o = n17106_o;
      7'b0000001: n17107_o = n17106_o;
      default: n17107_o = n17106_o;
    endcase
  assign n17108_o = dp_readdata_r[59:48];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17109_o = n17108_o;
      7'b0100000: n17109_o = n17108_o;
      7'b0010000: n17109_o = n17108_o;
      7'b0001000: n17109_o = n17086_o;
      7'b0000100: n17109_o = n17108_o;
      7'b0000010: n17109_o = n17108_o;
      7'b0000001: n17109_o = n17108_o;
      default: n17109_o = n17108_o;
    endcase
  assign n17110_o = dp_readdata_r[71:60];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17111_o = n17110_o;
      7'b0100000: n17111_o = n17110_o;
      7'b0010000: n17111_o = n17110_o;
      7'b0001000: n17111_o = n17110_o;
      7'b0000100: n17111_o = n17083_o;
      7'b0000010: n17111_o = n17110_o;
      7'b0000001: n17111_o = n17110_o;
      default: n17111_o = n17110_o;
    endcase
  assign n17112_o = dp_readdata_r[83:72];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17113_o = n17112_o;
      7'b0100000: n17113_o = n17112_o;
      7'b0010000: n17113_o = n17112_o;
      7'b0001000: n17113_o = n17112_o;
      7'b0000100: n17113_o = n17112_o;
      7'b0000010: n17113_o = n17080_o;
      7'b0000001: n17113_o = n17112_o;
      default: n17113_o = n17112_o;
    endcase
  assign n17114_o = dp_readdata_r[95:84];
  /* ../../HW/src/pcore/pcore.vhd:889:20  */
  always @*
    case (n17099_o)
      7'b1000000: n17115_o = n17114_o;
      7'b0100000: n17115_o = n17114_o;
      7'b0010000: n17115_o = n17114_o;
      7'b0001000: n17115_o = n17114_o;
      7'b0000100: n17115_o = n17114_o;
      7'b0000010: n17115_o = n17114_o;
      7'b0000001: n17115_o = n17077_o;
      default: n17115_o = n17114_o;
    endcase
  /* ../../HW/src/pcore/pcore.vhd:907:45  */
  assign n17117_o = dp_read_scatter_cnt_vm == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:907:20  */
  assign n17120_o = n17117_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n17121_o = dp_read_gen_valid_vm ? dp_readdata_vm : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:917:20  */
  assign n17122_o = dp_read_gen_valid_vm ? dp_readdata2_r : dp_readdata_vm;
  assign n17123_o = {n17115_o, n17113_o, n17111_o, n17109_o, n17107_o, n17105_o, n17103_o, n17101_o};
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n17124_o = n17075_o ? n17123_o : n17121_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n17125_o = n17075_o ? dp_readdata2_r : n17122_o;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n17127_o = n17075_o ? n17120_o : 1'b1;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n17129_o = n17075_o ? 3'b000 : dp_read_vector_vm;
  /* ../../HW/src/pcore/pcore.vhd:886:17  */
  assign n17131_o = n17075_o ? 3'b000 : dp_read_vaddr_vm;
  /* ../../HW/src/pcore/pcore.vhd:885:13  */
  assign n17136_o = dp_readena_vm ? n17127_o : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:958:26  */
  assign xregister_file_i_n17185 = xregister_file_i_read_result_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:959:24  */
  assign xregister_file_i_n17186 = xregister_file_i_read_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:945:1  */
  xregister_file xregister_file_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .write_result_vector_in(wr_vector),
    .write_result_lane_in(wr_vector_lane),
    .write_addr_in(result_write_addr),
    .write_result_ena_in(wr_flag1),
    .write_xreg_ena_in(wr_xreg1),
    .write_xreg_result_ena_in(wr_xreg_flag1),
    .write_data_in(mu_y),
    .write_result_in(mu_result),
    .read_addr_in(result_raddr1),
    .read_result_out(xregister_file_i_read_result_out),
    .read_xreg_out(xregister_file_i_read_xreg_out));
  /* ../../HW/src/pcore/pcore.vhd:975:27  */
  assign iregister_i_n17191 = iregister_i_rd_data1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:977:26  */
  assign iregister_i_n17192 = iregister_i_rd_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:967:1  */
  iregister_file iregister_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en1_in(i_rd_en1),
    .rd_vm_in(i_rd_vm),
    .rd_tid1_in(i_rd_tid1),
    .wr_tid1_in(i_wr_tid1),
    .wr_en1_in(i_wr_en1),
    .wr_vm_in(i_wr_vm),
    .wr_lane_in(wr_lane),
    .wr_addr1_in(i_wr_addr1),
    .wr_data1_in(i_wr_data1),
    .rd_data1_out(iregister_i_rd_data1_out),
    .rd_lane_out(iregister_i_rd_lane_out));
  /* ../../HW/src/pcore/pcore.vhd:993:14  */
  assign n17199_o = ~dp_rd_fork;
  /* ../../HW/src/pcore/pcore.vhd:994:33  */
  assign n17201_o = dp_rd_pid == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:994:20  */
  assign n17202_o = n17201_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:994:77  */
  assign n17204_o = dp_rd_cid == 3'b000;
  /* ../../HW/src/pcore/pcore.vhd:994:64  */
  assign n17205_o = n17204_o & n17202_o;
  /* ../../HW/src/pcore/pcore.vhd:994:4  */
  assign n17208_o = n17205_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1000:33  */
  assign n17210_o = dp_rd_pid == 2'b00;
  /* ../../HW/src/pcore/pcore.vhd:1000:20  */
  assign n17211_o = n17210_o & dp_read;
  /* ../../HW/src/pcore/pcore.vhd:1000:4  */
  assign n17214_o = n17211_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:993:1  */
  assign n17215_o = n17199_o ? n17208_o : n17214_o;
  /* ../../HW/src/pcore/pcore.vhd:1018:23  */
  assign n17223_o = dp_wr_mcast[4:0];
  /* ../../HW/src/pcore/pcore.vhd:1019:28  */
  assign n17224_o = dp_wr_mcast[5];
  /* ../../HW/src/pcore/pcore.vhd:1020:54  */
  assign n17225_o = dp_mcast_addr + n17223_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:36  */
  assign n17226_o = n17223_o & dp_mcast_addr;
  /* ../../HW/src/pcore/pcore.vhd:1030:64  */
  assign n17228_o = n17223_o & 5'b00000;
  /* ../../HW/src/pcore/pcore.vhd:1030:54  */
  assign n17229_o = n17226_o == n17228_o;
  /* ../../HW/src/pcore/pcore.vhd:1030:23  */
  assign n17230_o = n17229_o & n17224_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:18  */
  assign n17231_o = ~n17224_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:47  */
  assign n17233_o = $unsigned(5'b00000) >= $unsigned(dp_mcast_addr);
  /* ../../HW/src/pcore/pcore.vhd:1032:23  */
  assign n17234_o = n17233_o & n17231_o;
  /* ../../HW/src/pcore/pcore.vhd:1032:99  */
  assign n17236_o = $unsigned(5'b00000) <= $unsigned(n17225_o);
  /* ../../HW/src/pcore/pcore.vhd:1032:75  */
  assign n17237_o = n17236_o & n17234_o;
  /* ../../HW/src/pcore/pcore.vhd:1031:5  */
  assign n17238_o = n17230_o | n17237_o;
  /* ../../HW/src/pcore/pcore.vhd:1028:20  */
  assign n17239_o = n17238_o & dp_write;
  /* ../../HW/src/pcore/pcore.vhd:1028:1  */
  assign n17242_o = n17239_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/pcore.vhd:1050:51  */
  assign n17245_o = xreg_read[31:0];
  /* ../../HW/src/pcore/pcore.vhd:1051:45  */
  assign n17246_o = mu_x1[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1052:45  */
  assign n17247_o = mu_x2[11:0];
  /* ../../HW/src/pcore/pcore.vhd:1054:40  */
  assign alu_0_i_n17248 = alu_0_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1055:41  */
  assign alu_0_i_n17249 = alu_0_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1056:41  */
  assign alu_0_i_n17250 = alu_0_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1046:1  */
  alu alu_0_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17245_o),
    .x1_in(n17246_o),
    .x2_in(n17247_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_0_i_y_out),
    .y2_out(alu_0_i_y2_out),
    .y3_out(alu_0_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1062:51  */
  assign n17257_o = xreg_read[63:32];
  /* ../../HW/src/pcore/pcore.vhd:1063:45  */
  assign n17258_o = mu_x1[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1064:45  */
  assign n17259_o = mu_x2[23:12];
  /* ../../HW/src/pcore/pcore.vhd:1066:40  */
  assign alu_1_i_n17260 = alu_1_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1067:41  */
  assign alu_1_i_n17261 = alu_1_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1068:41  */
  assign alu_1_i_n17262 = alu_1_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1058:1  */
  alu alu_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17257_o),
    .x1_in(n17258_o),
    .x2_in(n17259_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_1_i_y_out),
    .y2_out(alu_1_i_y2_out),
    .y3_out(alu_1_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1074:51  */
  assign n17269_o = xreg_read[95:64];
  /* ../../HW/src/pcore/pcore.vhd:1075:45  */
  assign n17270_o = mu_x1[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1076:45  */
  assign n17271_o = mu_x2[35:24];
  /* ../../HW/src/pcore/pcore.vhd:1078:40  */
  assign alu_2_i_n17272 = alu_2_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1079:41  */
  assign alu_2_i_n17273 = alu_2_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1080:41  */
  assign alu_2_i_n17274 = alu_2_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1070:1  */
  alu alu_2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17269_o),
    .x1_in(n17270_o),
    .x2_in(n17271_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_2_i_y_out),
    .y2_out(alu_2_i_y2_out),
    .y3_out(alu_2_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1086:51  */
  assign n17281_o = xreg_read[127:96];
  /* ../../HW/src/pcore/pcore.vhd:1087:45  */
  assign n17282_o = mu_x1[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1088:45  */
  assign n17283_o = mu_x2[47:36];
  /* ../../HW/src/pcore/pcore.vhd:1090:40  */
  assign alu_3_i_n17284 = alu_3_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1091:41  */
  assign alu_3_i_n17285 = alu_3_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1092:41  */
  assign alu_3_i_n17286 = alu_3_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1082:1  */
  alu alu_3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17281_o),
    .x1_in(n17282_o),
    .x2_in(n17283_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_3_i_y_out),
    .y2_out(alu_3_i_y2_out),
    .y3_out(alu_3_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1098:51  */
  assign n17293_o = xreg_read[159:128];
  /* ../../HW/src/pcore/pcore.vhd:1099:45  */
  assign n17294_o = mu_x1[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1100:45  */
  assign n17295_o = mu_x2[59:48];
  /* ../../HW/src/pcore/pcore.vhd:1102:40  */
  assign alu_4_i_n17296 = alu_4_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1103:41  */
  assign alu_4_i_n17297 = alu_4_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1104:41  */
  assign alu_4_i_n17298 = alu_4_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1094:1  */
  alu alu_4_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17293_o),
    .x1_in(n17294_o),
    .x2_in(n17295_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_4_i_y_out),
    .y2_out(alu_4_i_y2_out),
    .y3_out(alu_4_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1110:51  */
  assign n17305_o = xreg_read[191:160];
  /* ../../HW/src/pcore/pcore.vhd:1111:45  */
  assign n17306_o = mu_x1[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1112:45  */
  assign n17307_o = mu_x2[71:60];
  /* ../../HW/src/pcore/pcore.vhd:1114:40  */
  assign alu_5_i_n17308 = alu_5_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1115:41  */
  assign alu_5_i_n17309 = alu_5_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1116:41  */
  assign alu_5_i_n17310 = alu_5_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1106:1  */
  alu alu_5_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17305_o),
    .x1_in(n17306_o),
    .x2_in(n17307_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_5_i_y_out),
    .y2_out(alu_5_i_y2_out),
    .y3_out(alu_5_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1122:51  */
  assign n17317_o = xreg_read[223:192];
  /* ../../HW/src/pcore/pcore.vhd:1123:45  */
  assign n17318_o = mu_x1[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1124:45  */
  assign n17319_o = mu_x2[83:72];
  /* ../../HW/src/pcore/pcore.vhd:1126:40  */
  assign alu_6_i_n17320 = alu_6_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1127:41  */
  assign alu_6_i_n17321 = alu_6_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1128:41  */
  assign alu_6_i_n17322 = alu_6_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1118:1  */
  alu alu_6_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17317_o),
    .x1_in(n17318_o),
    .x2_in(n17319_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_6_i_y_out),
    .y2_out(alu_6_i_y2_out),
    .y3_out(alu_6_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1134:51  */
  assign n17329_o = xreg_read[255:224];
  /* ../../HW/src/pcore/pcore.vhd:1135:45  */
  assign n17330_o = mu_x1[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1136:45  */
  assign n17331_o = mu_x2[95:84];
  /* ../../HW/src/pcore/pcore.vhd:1138:40  */
  assign alu_7_i_n17332 = alu_7_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1139:41  */
  assign alu_7_i_n17333 = alu_7_i_y2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1140:41  */
  assign alu_7_i_n17334 = alu_7_i_y3_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1130:1  */
  alu alu_7_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .mu_opcode_in(mu_opcodes),
    .mu_tid_in(mu_tid),
    .xreg_in(n17329_o),
    .x1_in(n17330_o),
    .x2_in(n17331_o),
    .x_scalar_in(mu_x_scalar),
    .y_out(alu_7_i_y_out),
    .y2_out(alu_7_i_y2_out),
    .y3_out(alu_7_i_y3_out));
  /* ../../HW/src/pcore/pcore.vhd:1143:24  */
  assign n17341_o = i_y_neg & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1145:26  */
  assign n17342_o = i_y_zero & enable_in;
  /* ../../HW/src/pcore/pcore.vhd:1156:34  */
  assign ialu_i_n17343 = ialu_i_y_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1157:38  */
  assign ialu_i_n17344 = ialu_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1158:39  */
  assign ialu_i_n17345 = ialu_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1151:1  */
  ialu ialu_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(i_opcode),
    .x1_in(i_x1),
    .x2_in(i_x2),
    .y_out(ialu_i_y_out),
    .y_neg_out(ialu_i_y_neg_out),
    .y_zero_out(ialu_i_y_zero_out));
  /* ../../HW/src/pcore/pcore.vhd:1182:27  */
  assign register_bank_i_n17354 = register_bank_i_rd_x1_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1183:27  */
  assign register_bank_i_n17355 = register_bank_i_rd_x2_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1201:39  */
  assign n17356_o = gen_rd_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1203:39  */
  assign n17357_o = gen_wr_addr_r[16:0];
  /* ../../HW/src/pcore/pcore.vhd:1209:28  */
  assign register_bank_i_n17358 = register_bank_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1210:31  */
  assign register_bank_i_n17359 = register_bank_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1211:27  */
  assign register_bank_i_n17360 = register_bank_i_dp_readena_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1212:31  */
  assign register_bank_i_n17361 = register_bank_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1213:30  */
  assign register_bank_i_n17362 = register_bank_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1214:32  */
  assign register_bank_i_n17363 = register_bank_i_dp_read_scatter_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1215:36  */
  assign register_bank_i_n17364 = register_bank_i_dp_read_scatter_cnt_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1216:39  */
  assign register_bank_i_n17365 = register_bank_i_dp_read_scatter_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1217:34  */
  assign register_bank_i_n17366 = register_bank_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1218:34  */
  assign register_bank_i_n17367 = register_bank_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1219:34  */
  assign register_bank_i_n17368 = register_bank_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1220:31  */
  assign register_bank_i_n17369 = register_bank_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1221:34  */
  assign register_bank_i_n17370 = register_bank_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1169:1  */
  register_bank register_bank_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .rd_en_in(rd_en1),
    .rd_en_vm_in(rd_vm),
    .rd_x1_vector_in(rd_x1_vector1),
    .rd_x1_addr_in(rd_x1_addr1),
    .rd_x2_vector_in(rd_x2_vector1),
    .rd_x2_addr_in(rd_x2_addr1),
    .wr_en_in(wr_en1),
    .wr_en_vm_in(wr_vm),
    .wr_vector_in(wr_vector),
    .wr_addr_in(wr_addr1),
    .wr_data_in(wr_data1),
    .wr_lane_in(wr_vector_lane),
    .dp_rd_vector_in(gen_read_vector_r),
    .dp_rd_scatter_in(gen_read_scatter_r),
    .dp_rd_scatter_cnt_in(gen_read_scatter_cnt_r),
    .dp_rd_scatter_vector_in(gen_read_scatter_vector_r),
    .dp_rd_gen_valid_in(gen_read_gen_valid_r),
    .dp_rd_data_flow_in(gen_read_data_flow_r),
    .dp_rd_data_type_in(gen_read_data_type_r),
    .dp_rd_stream_in(gen_read_stream_r),
    .dp_rd_stream_id_in(gen_read_stream_id_r),
    .dp_rd_addr_in(n17356_o),
    .dp_wr_vector_in(gen_write_vector_r),
    .dp_wr_addr_in(n17357_o),
    .dp_write_in(gen_write_r),
    .dp_write_vm_in(gen_write_vm_r),
    .dp_read_in(gen_read_r),
    .dp_read_vm_in(gen_read_vm_r),
    .dp_writedata_in(gen_writedata_r),
    .rd_en_out(),
    .rd_x1_data_out(register_bank_i_rd_x1_data_out),
    .rd_x2_data_out(register_bank_i_rd_x2_data_out),
    .dp_readdata_out(register_bank_i_dp_readdata_out),
    .dp_readdata_vm_out(register_bank_i_dp_readdata_vm_out),
    .dp_readena_out(register_bank_i_dp_readena_out),
    .dp_read_vector_out(register_bank_i_dp_read_vector_out),
    .dp_read_vaddr_out(register_bank_i_dp_read_vaddr_out),
    .dp_read_scatter_out(register_bank_i_dp_read_scatter_out),
    .dp_read_scatter_cnt_out(register_bank_i_dp_read_scatter_cnt_out),
    .dp_read_scatter_vector_out(register_bank_i_dp_read_scatter_vector_out),
    .dp_read_gen_valid_out(register_bank_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(register_bank_i_dp_read_data_flow_out),
    .dp_read_data_type_out(register_bank_i_dp_read_data_type_out),
    .dp_read_stream_out(register_bank_i_dp_read_stream_out),
    .dp_read_stream_id_out(register_bank_i_dp_read_stream_id_out));
  /* ../../HW/src/pcore/pcore.vhd:1253:60  */
  assign instr_decoder2_i_n17403 = instr_decoder2_i_opcode1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1254:56  */
  assign instr_decoder2_i_n17404 = instr_decoder2_i_en1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1256:68  */
  assign instr_decoder2_i_n17405 = instr_decoder2_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1257:58  */
  assign instr_decoder2_i_n17406 = instr_decoder2_i_xreg1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1258:58  */
  assign instr_decoder2_i_n17407 = instr_decoder2_i_flag1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1259:57  */
  assign instr_decoder2_i_n17408 = instr_decoder2_i_wren_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1261:55  */
  assign instr_decoder2_i_n17409 = instr_decoder2_i_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1263:61  */
  assign instr_decoder2_i_n17410 = instr_decoder2_i_x1_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1264:61  */
  assign instr_decoder2_i_n17411 = instr_decoder2_i_x2_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1265:60  */
  assign instr_decoder2_i_n17412 = instr_decoder2_i_y_addr1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1267:62  */
  assign instr_decoder2_i_n17413 = instr_decoder2_i_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1268:62  */
  assign instr_decoder2_i_n17414 = instr_decoder2_i_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1269:61  */
  assign instr_decoder2_i_n17415 = instr_decoder2_i_y_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1270:64  */
  assign instr_decoder2_i_n17416 = instr_decoder2_i_vector_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1273:61  */
  assign instr_decoder2_i_n17417 = instr_decoder2_i_x1_c1_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1274:58  */
  assign instr_decoder2_i_n17418 = instr_decoder2_i_x1_c1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1277:60  */
  assign instr_decoder2_i_n17419 = instr_decoder2_i_i_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1278:60  */
  assign instr_decoder2_i_n17420 = instr_decoder2_i_i_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1279:61  */
  assign instr_decoder2_i_n17421 = instr_decoder2_i_i_rd_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1281:61  */
  assign instr_decoder2_i_n17422 = instr_decoder2_i_i_wr_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1282:60  */
  assign instr_decoder2_i_n17423 = instr_decoder2_i_i_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1283:60  */
  assign instr_decoder2_i_n17424 = instr_decoder2_i_i_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1284:62  */
  assign instr_decoder2_i_n17425 = instr_decoder2_i_i_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1285:62  */
  assign instr_decoder2_i_n17426 = instr_decoder2_i_i_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1289:60  */
  assign instr_decoder2_i_n17427 = instr_decoder2_i_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1292:61  */
  assign instr_decoder2_i_n17428 = instr_decoder2_i_i_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1293:57  */
  assign instr_decoder2_i_n17429 = instr_decoder2_i_i_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1294:57  */
  assign instr_decoder2_i_n17430 = instr_decoder2_i_i_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1299:65  */
  assign instr_decoder2_i_n17431 = instr_decoder2_i_result_raddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1298:65  */
  assign instr_decoder2_i_n17432 = instr_decoder2_i_result_waddr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1230:1  */
  instr_decoder2_0_0 instr_decoder2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_r),
    .instruction_imu_in(instruction_imu_r),
    .instruction_mu_valid_in(instruction_mu_valid_r),
    .instruction_imu_valid_in(instruction_imu_valid_r),
    .instruction_tid_in(tid_r),
    .instruction_tid_valid_in(tid_valid1),
    .instruction_vm_in(vm_r),
    .instruction_data_model_in(data_model_r),
    .instruction_pre_pre_vm_in(pre_pre_vm_r),
    .instruction_pre_pre_data_model_in(pre_pre_data_model_r),
    .instruction_pre_tid_in(pre_tid_r),
    .instruction_pre_tid_valid_in(pre_tid_valid1),
    .instruction_pre_pre_tid_in(pre_pre_tid_r),
    .instruction_pre_pre_tid_valid_in(pre_pre_tid_valid1),
    .instruction_pre_iregister_auto_in(pre_iregister_auto_r),
    .i_rd_data_in(i_rd_data1),
    .lane_in(rd_lane),
    .i_y_in(i_y),
    .result_in(result_read),
    .opcode1_out(instr_decoder2_i_opcode1_out),
    .en1_out(instr_decoder2_i_en1_out),
    .instruction_tid_out(instr_decoder2_i_instruction_tid_out),
    .xreg1_out(instr_decoder2_i_xreg1_out),
    .flag1_out(instr_decoder2_i_flag1_out),
    .wren_out(instr_decoder2_i_wren_out),
    .vm_out(instr_decoder2_i_vm_out),
    .x1_addr1_out(instr_decoder2_i_x1_addr1_out),
    .x2_addr1_out(instr_decoder2_i_x2_addr1_out),
    .y_addr1_out(instr_decoder2_i_y_addr1_out),
    .x1_vector_out(instr_decoder2_i_x1_vector_out),
    .x2_vector_out(instr_decoder2_i_x2_vector_out),
    .y_vector_out(instr_decoder2_i_y_vector_out),
    .vector_lane_out(instr_decoder2_i_vector_lane_out),
    .x1_c1_en_out(instr_decoder2_i_x1_c1_en_out),
    .x1_c1_out(instr_decoder2_i_x1_c1_out),
    .i_rd_en_out(instr_decoder2_i_i_rd_en_out),
    .i_rd_vm_out(instr_decoder2_i_i_rd_vm_out),
    .i_rd_tid_out(instr_decoder2_i_i_rd_tid_out),
    .i_wr_tid_out(instr_decoder2_i_i_wr_tid_out),
    .i_wr_en_out(instr_decoder2_i_i_wr_en_out),
    .i_wr_vm_out(instr_decoder2_i_i_wr_vm_out),
    .i_wr_addr_out(instr_decoder2_i_i_wr_addr_out),
    .i_wr_data_out(instr_decoder2_i_i_wr_data_out),
    .wr_lane_out(instr_decoder2_i_wr_lane_out),
    .i_opcode_out(instr_decoder2_i_i_opcode_out),
    .i_x1_out(instr_decoder2_i_i_x1_out),
    .i_x2_out(instr_decoder2_i_i_x2_out),
    .result_waddr_out(instr_decoder2_i_result_waddr_out),
    .result_raddr_out(instr_decoder2_i_result_raddr_out));
  /* ../../HW/src/pcore/pcore.vhd:1332:26  */
  assign instr_dispatch2_i1_n17493 = instr_dispatch2_i1_rd_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1333:26  */
  assign instr_dispatch2_i1_n17494 = instr_dispatch2_i1_rd_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1334:31  */
  assign instr_dispatch2_i1_n17495 = instr_dispatch2_i1_rd_x1_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1335:31  */
  assign instr_dispatch2_i1_n17496 = instr_dispatch2_i1_rd_x2_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1339:33  */
  assign instr_dispatch2_i1_n17497 = instr_dispatch2_i1_rd_x1_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1340:33  */
  assign instr_dispatch2_i1_n17498 = instr_dispatch2_i1_rd_x2_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1347:28  */
  assign instr_dispatch2_i1_n17499 = instr_dispatch2_i1_wr_xreg_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1348:28  */
  assign instr_dispatch2_i1_n17500 = instr_dispatch2_i1_wr_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1349:33  */
  assign instr_dispatch2_i1_n17501 = instr_dispatch2_i1_wr_xreg_flag_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1350:26  */
  assign instr_dispatch2_i1_n17502 = instr_dispatch2_i1_wr_en_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1351:26  */
  assign instr_dispatch2_i1_n17503 = instr_dispatch2_i1_wr_vm_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1352:30  */
  assign instr_dispatch2_i1_n17504 = instr_dispatch2_i1_wr_vector_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1353:28  */
  assign instr_dispatch2_i1_n17505 = instr_dispatch2_i1_wr_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1354:35  */
  assign instr_dispatch2_i1_n17506 = instr_dispatch2_i1_wr_result_addr_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1355:28  */
  assign instr_dispatch2_i1_n17507 = instr_dispatch2_i1_wr_data_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1356:28  */
  assign instr_dispatch2_i1_n17508 = instr_dispatch2_i1_wr_lane_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1358:26  */
  assign instr_dispatch2_i1_n17509 = instr_dispatch2_i1_mu_x1_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1359:26  */
  assign instr_dispatch2_i1_n17510 = instr_dispatch2_i1_mu_x2_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1360:32  */
  assign instr_dispatch2_i1_n17511 = instr_dispatch2_i1_mu_x_scalar_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1361:30  */
  assign instr_dispatch2_i1_n17512 = instr_dispatch2_i1_mu_opcode_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1362:27  */
  assign instr_dispatch2_i1_n17513 = instr_dispatch2_i1_mu_tid_out; // (signal)
  /* ../../HW/src/pcore/pcore.vhd:1309:1  */
  instr_dispatch2 instr_dispatch2_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .opcode_in(opcode1),
    .instruction_tid_in(tid_decoder2dispatch),
    .xreg_in(mu_xreg1),
    .flag_in(mu_flag1),
    .wren_in(mu_wren),
    .en_in(en1),
    .vm_in(mu_vm),
    .x1_addr1_in(x1_addr1),
    .x2_addr1_in(x2_addr1),
    .y_addr1_in(y_addr1),
    .result_addr1_in(result_waddr1),
    .x1_vector_in(x1_vector),
    .x2_vector_in(x2_vector),
    .y_vector_in(y_vector),
    .vector_lane_in(vector_lane),
    .x1_c1_en_in(x1_c1_en),
    .x1_c1_in(x1_c1),
    .rd_x1_data_in(rd_x1_data1),
    .rd_x2_data_in(rd_x2_data1),
    .mu_y_in(mu_y2),
    .rd_en_out(instr_dispatch2_i1_rd_en_out),
    .rd_vm_out(instr_dispatch2_i1_rd_vm_out),
    .rd_x1_addr_out(instr_dispatch2_i1_rd_x1_addr_out),
    .rd_x2_addr_out(instr_dispatch2_i1_rd_x2_addr_out),
    .rd_x1_vector_out(instr_dispatch2_i1_rd_x1_vector_out),
    .rd_x2_vector_out(instr_dispatch2_i1_rd_x2_vector_out),
    .wr_xreg_out(instr_dispatch2_i1_wr_xreg_out),
    .wr_flag_out(instr_dispatch2_i1_wr_flag_out),
    .wr_xreg_flag_out(instr_dispatch2_i1_wr_xreg_flag_out),
    .wr_en_out(instr_dispatch2_i1_wr_en_out),
    .wr_vm_out(instr_dispatch2_i1_wr_vm_out),
    .wr_vector_out(instr_dispatch2_i1_wr_vector_out),
    .wr_addr_out(instr_dispatch2_i1_wr_addr_out),
    .wr_result_addr_out(instr_dispatch2_i1_wr_result_addr_out),
    .wr_data_out(instr_dispatch2_i1_wr_data_out),
    .wr_lane_out(instr_dispatch2_i1_wr_lane_out),
    .mu_x1_out(instr_dispatch2_i1_mu_x1_out),
    .mu_x2_out(instr_dispatch2_i1_mu_x2_out),
    .mu_x_scalar_out(instr_dispatch2_i1_mu_x_scalar_out),
    .mu_opcode_out(instr_dispatch2_i1_mu_opcode_out),
    .mu_tid_out(instr_dispatch2_i1_mu_tid_out));
  assign n17559_o = {alu_7_i_n17332, alu_6_i_n17320, alu_5_i_n17308, alu_4_i_n17296, alu_3_i_n17284, alu_2_i_n17272, alu_1_i_n17260, alu_0_i_n17248};
  assign n17560_o = {alu_7_i_n17334, alu_6_i_n17322, alu_5_i_n17310, alu_4_i_n17298, alu_3_i_n17286, alu_2_i_n17274, alu_1_i_n17262, alu_0_i_n17250};
  assign n17561_o = {alu_7_i_n17333, alu_6_i_n17321, alu_5_i_n17309, alu_4_i_n17297, alu_3_i_n17285, alu_2_i_n17273, alu_1_i_n17261, alu_0_i_n17249};
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17562_o = dp_readena_vm ? n17124_o : dp_readdata_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17563_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n17563_q <= n17562_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17564_o = dp_readena_vm ? n17125_o : dp_readdata2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17565_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n17565_q <= n17564_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17566_q <= 1'b0;
    else
      n17566_q <= n17136_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17567_q <= 1'b0;
    else
      n17567_q <= dp_readdata_vm_vm;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17568_o = dp_readena_vm ? dp_read_gen_valid_vm : dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17569_q <= 1'b0;
    else
      n17569_q <= n17568_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17570_o = dp_readena_vm ? dp_read_data_flow_vm : dp_read_data_flow2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17571_q <= 2'b00;
    else
      n17571_q <= n17570_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17572_o = dp_readena_vm ? dp_read_data_type_vm : dp_read_data_type2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17573_q <= 2'b00;
    else
      n17573_q <= n17572_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17574_o = dp_readena_vm ? n17129_o : dp_read_vector2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17575_q <= 3'b000;
    else
      n17575_q <= n17574_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17576_o = dp_readena_vm ? n17131_o : dp_read_vaddr2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17577_q <= 3'b000;
    else
      n17577_q <= n17576_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17578_o = dp_readena_vm ? dp_read_stream_vm : dp_read_stream2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17579_q <= 1'b0;
    else
      n17579_q <= n17578_o;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  assign n17580_o = dp_readena_vm ? dp_read_stream_id_vm : dp_read_stream_id2_r;
  /* ../../HW/src/pcore/pcore.vhd:883:9  */
  always @(posedge clock_in or posedge n17072_o)
    if (n17072_o)
      n17581_q <= 2'b00;
    else
      n17581_q <= n17580_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17582_q <= 3'b000;
    else
      n17582_q <= write_scatter_curr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17583_q <= 3'b000;
    else
      n17583_q <= dp_read_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17584_q <= 2'b00;
    else
      n17584_q <= dp_read_scatter;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17587_q <= 3'b000;
    else
      n17587_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17588_q <= 3'b000;
    else
      n17588_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17589_q <= 1'b0;
    else
      n17589_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17590_q <= 2'b00;
    else
      n17590_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17591_q <= 2'b00;
    else
      n17591_q <= dp_read_data_type;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17592_q <= 1'b0;
    else
      n17592_q <= dp_read_stream;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17593_q <= 2'b00;
    else
      n17593_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17594_q <= 22'b0000000000000000000000;
    else
      n17594_q <= dp_rd_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17595_q <= 3'b000;
    else
      n17595_q <= dp_write_vector;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17596_q <= 22'b0000000000000000000000;
    else
      n17596_q <= dp_wr_addr;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17597_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n17597_q <= dp_writedata;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17598_o = n16745_o ? dp_rd_vm : dp_rd_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17599_q <= 1'b0;
    else
      n17599_q <= n17598_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17600_o = n16745_o ? dp_rd_fork : dp_rd_fork_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17601_q <= 1'b0;
    else
      n17601_q <= n17600_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17602_o = n16891_o ? dp_wr_vm : dp_wr_vm_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17603_q <= 1'b0;
    else
      n17603_q <= n17602_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17606_q <= 22'b0000000000000000000000;
    else
      n17606_q <= n16743_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17607_q <= 22'b0000000000000000000000;
    else
      n17607_q <= n16889_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17608_o = n16891_o ? dp_wr_mcast : dp_wr_mcast_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17609_q <= 6'b000000;
    else
      n17609_q <= n17608_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17610_o = n16891_o ? dp_write : dp_write_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17611_q <= 1'b0;
    else
      n17611_q <= n17610_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17614_o = n16891_o ? dp_write_vector : dp_write_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17615_q <= 3'b000;
    else
      n17615_q <= n17614_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17616_o = n16891_o ? dp_write_scatter : dp_write_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17617_q <= 2'b00;
    else
      n17617_q <= n17616_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17618_o = n16891_o ? dp_write_share : dp_write_share_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17619_q <= 1'b0;
    else
      n17619_q <= n17618_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  assign n17620_o = n16891_o ? dp_write_step : dp_write_step_r;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17621_q <= 22'b0000000000000000000000;
    else
      n17621_q <= n17620_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17622_o = n16745_o ? dp_read : dp_read_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17623_q <= 1'b0;
    else
      n17623_q <= n17622_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17624_o = n16745_o ? dp_read_vector : dp_read_vector_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17625_q <= 3'b000;
    else
      n17625_q <= n17624_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17626_o = n16745_o ? dp_read_scatter : dp_read_scatter_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17627_q <= 2'b00;
    else
      n17627_q <= n17626_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n17628_o = ~n16732_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n17629_o = n16745_o & n17628_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17630_o = n17629_o ? dp_read_share : dp_read_share_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n17631_q <= n17630_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n17632_o = ~n16732_o;
  /* ../../HW/src/pcore/pcore.vhd:570:1  */
  assign n17633_o = n16745_o & n17632_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17634_o = n17633_o ? dp_read_step : dp_read_step_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in)
    n17635_q <= n17634_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17636_o = n16745_o ? dp_read_gen_valid : dp_read_gen_valid_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17637_q <= 1'b0;
    else
      n17637_q <= n17636_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17638_o = n16745_o ? dp_read_data_flow : dp_read_data_flow_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17639_q <= 2'b00;
    else
      n17639_q <= n17638_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17640_o = n16745_o ? dp_read_data_type : dp_read_data_type_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17641_q <= 2'b00;
    else
      n17641_q <= n17640_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17642_o = n16745_o ? dp_read_stream : dp_read_stream_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17643_q <= 1'b0;
    else
      n17643_q <= n17642_o;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  assign n17644_o = n16745_o ? dp_read_stream_id : dp_read_stream_id_r;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17645_q <= 2'b00;
    else
      n17645_q <= n17644_o;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17646_q <= 84'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n17646_q <= n16903_o;
  /* ../../HW/src/pcore/pcore.vhd:690:4  */
  assign n17647_o = {n16946_o, n17646_q};
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17648_q <= 3'b000;
    else
      n17648_q <= read_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:588:7  */
  always @(posedge clock_in or posedge n16732_o)
    if (n16732_o)
      n17649_q <= 3'b000;
    else
      n17649_q <= read_scatter_vector;
  /* ../../HW/src/pcore/pcore.vhd:706:7  */
  always @(posedge clock_in or posedge n16878_o)
    if (n16878_o)
      n17650_q <= 3'b000;
    else
      n17650_q <= write_scatter_cnt;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17652_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n17652_q <= instruction_mu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17653_q <= 32'b00000000000000000000000000000000;
    else
      n17653_q <= instruction_imu_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17654_q <= 1'b0;
    else
      n17654_q <= instruction_mu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17655_q <= 1'b0;
    else
      n17655_q <= instruction_imu_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17656_q <= 1'b0;
    else
      n17656_q <= vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17657_q <= 2'b00;
    else
      n17657_q <= data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17658_q <= 4'b0000;
    else
      n17658_q <= tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17659_q <= 1'b0;
    else
      n17659_q <= tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17660_q <= 4'b0000;
    else
      n17660_q <= pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17661_q <= 1'b0;
    else
      n17661_q <= pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17662_q <= 4'b0000;
    else
      n17662_q <= pre_pre_tid_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17663_q <= 1'b0;
    else
      n17663_q <= pre_pre_tid_valid1_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17664_q <= 1'b0;
    else
      n17664_q <= pre_pre_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17665_q <= 2'b00;
    else
      n17665_q <= pre_pre_data_model_in;
  /* ../../HW/src/pcore/pcore.vhd:842:9  */
  always @(posedge clock_in or posedge n17021_o)
    if (n17021_o)
      n17666_q <= 28'b0000000000000000000000000000;
    else
      n17666_q <= pre_iregister_auto_in;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17667_q <= 1'b0;
    else
      n17667_q <= write;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17668_q <= 1'b0;
    else
      n17668_q <= dp_wr_vm;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17670_q <= 1'b0;
    else
      n17670_q <= read;
  /* ../../HW/src/pcore/pcore.vhd:653:7  */
  always @(posedge clock_in or posedge n16809_o)
    if (n16809_o)
      n17671_q <= 1'b0;
    else
      n17671_q <= dp_rd_vm;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17673_q <= 1'b0;
    else
      n17673_q <= dp_rd_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17674_q <= 1'b0;
    else
      n17674_q <= dp_wr_vm_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17675_q <= 1'b0;
    else
      n17675_q <= dp_code_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17676_q <= 22'b0000000000000000000000;
    else
      n17676_q <= dp_rd_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17677_q <= 1'b0;
    else
      n17677_q <= dp_rd_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17678_q <= 22'b0000000000000000000000;
    else
      n17678_q <= dp_rd_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17679_q <= 22'b0000000000000000000000;
    else
      n17679_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17680_q <= 1'b0;
    else
      n17680_q <= dp_wr_share_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17681_q <= 22'b0000000000000000000000;
    else
      n17681_q <= dp_wr_addr_step_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17682_q <= 6'b000000;
    else
      n17682_q <= dp_wr_mcast_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17683_q <= 1'b0;
    else
      n17683_q <= dp_write_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17684_q <= 1'b0;
    else
      n17684_q <= dp_wr_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17685_q <= 1'b0;
    else
      n17685_q <= dp_write_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17686_q <= 3'b000;
    else
      n17686_q <= dp_write_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17687_q <= 2'b00;
    else
      n17687_q <= dp_write_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17688_q <= 1'b0;
    else
      n17688_q <= dp_rd_fork_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17689_q <= 1'b0;
    else
      n17689_q <= dp_read_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17690_q <= 3'b000;
    else
      n17690_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17691_q <= 2'b00;
    else
      n17691_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17692_q <= 1'b0;
    else
      n17692_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17693_q <= 2'b00;
    else
      n17693_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17694_q <= 2'b00;
    else
      n17694_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17695_q <= 1'b0;
    else
      n17695_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17696_q <= 2'b00;
    else
      n17696_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17697_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n17697_q <= dp_writedata_in;
  /* ../../HW/src/pcore/pcore.vhd:377:4  */
  always @(posedge clock_in or posedge n16536_o)
    if (n16536_o)
      n17698_q <= 1'b0;
    else
      n17698_q <= dp_config_in_in;
  /* ../../HW/src/pcore/pcore.vhd:796:41  */
  assign n17699_o = dp_readena_r ? dp_read_vector2_r : 3'bz;
  /* ../../HW/src/pcore/pcore.vhd:797:39  */
  assign n17700_o = dp_readena_r ? dp_read_vaddr2_r : 3'bz;
endmodule

module instr_fetch
  (input  clock_in,
   input  reset_in,
   input  [127:0] rom_data_in,
   input  [10:0] task_start_addr_in,
   input  task_in,
   input  [4:0] task_pcore_max_in,
   input  task_vm_in,
   input  task_lockstep_in,
   input  [3:0] task_tid_mask_in,
   input  [27:0] task_iregister_auto_in,
   input  [1:0] task_data_model_in,
   input  i_y_neg_in,
   input  i_y_zero_in,
   output [79:0] instruction_mu_out,
   output [31:0] instruction_imu_out,
   output instruction_mu_valid_out,
   output instruction_imu_valid_out,
   output instruction_vm_out,
   output [1:0] instruction_data_model_out,
   output [3:0] instruction_tid_out,
   output instruction_tid_valid_out,
   output [3:0] instruction_pre_tid_out,
   output instruction_pre_tid_valid_out,
   output [3:0] instruction_pre_pre_tid_out,
   output instruction_pre_pre_tid_valid_out,
   output instruction_pre_pre_vm_out,
   output [1:0] instruction_pre_pre_data_model_out,
   output [7:0] instruction_pcore_enable_out,
   output [27:0] instruction_pre_iregister_auto_out,
   output [10:0] rom_addr_out,
   output [10:0] rom_addr_plus_2_out,
   output [1:0] busy_out,
   output ready_out);
  wire [175:0] pc_r;
  wire [15:0] busy_r;
  wire [15:0] vm_r;
  wire [15:0] vm_rr;
  wire [31:0] data_model_r;
  wire [31:0] data_model_rr;
  wire [447:0] iregister_auto_r;
  wire [447:0] iregister_auto_rr;
  wire [15:0] tid;
  wire [15:0] tid_delay;
  wire [15:0] tid_r;
  wire tid_valid_r;
  wire [15:0] tid_rr;
  wire tid_valid_rr;
  wire tid_valid_rrr;
  wire [15:0] tid_rrr;
  wire [15:0] tid_rrrr;
  wire [15:0] tid_rrrrr;
  wire [15:0] tid_rrrrrr;
  wire [15:0] tid_rrrrrrr;
  wire [15:0] tid_rrrrrrrr;
  wire [15:0] tid_rrrrrrrrr;
  wire [15:0] tid_rrrrrrrrrr;
  wire [15:0] tid_rrrrrrrrrrr;
  wire [3:0] tid2_r;
  wire [3:0] tid2_rr;
  wire [3:0] tid2_rrr;
  wire [10:0] rom_addr;
  wire [10:0] rom_addr_r;
  wire [10:0] rom_addr_rr;
  wire [15:0] delay_r;
  wire [15:0] busy1;
  wire [1:0] busy2;
  wire [1:0] busy2_r;
  wire [15:0] avail;
  wire [15:0] avail_r;
  wire [15:0] next_tid;
  wire [3:0] next_tid2;
  wire next_tid_valid;
  wire [79:0] instruction_mu_r;
  wire [31:0] instruction_imu_r;
  wire instruction_mu_valid_r;
  wire instruction_imu_valid_r;
  wire [10:0] task_start_addr_r;
  wire [4:0] task_pcore_max_r;
  wire [4:0] task_pcore_curr_r;
  reg [15:0] task_tid_mask_r;
  wire [15:0] task_tid_mask;
  wire task_lockstep_r;
  wire [15:0] task_mask_r;
  wire task_vm_r;
  wire [27:0] task_iregister_auto_r;
  wire [1:0] task2_data_model_r;
  wire [79:0] mu_instruction;
  wire [31:0] imu_instruction;
  wire [15:0] ctrl_instruction;
  wire [10:0] instruction_addr_r;
  wire [10:0] instruction_addr_rr;
  wire got_control_r;
  wire got_control_rr;
  wire got_control_rrr;
  wire got_control_rrrr;
  wire got_control_rrrrr;
  wire got_control_rrrrrr;
  wire got_control_rrrrrrr;
  wire got_control_rrrrrrrr;
  wire [4:0] ctrl_opcode_r;
  wire [10:0] ctrl_goto_addr_r;
  wire [4:0] ctrl_opcode_rr;
  wire [10:0] ctrl_goto_addr_rr;
  wire [4:0] ctrl_opcode_rrr;
  wire [10:0] ctrl_goto_addr_rrr;
  wire [10:0] ctrl_next_addr_r;
  wire [10:0] ctrl_next_addr_rr;
  wire [10:0] ctrl_next_addr_rrr;
  wire [10:0] ctrl_next_addr_rrrr;
  wire [10:0] ctrl_next_addr_rrrrr;
  wire [10:0] ctrl_next_addr_rrrrrr;
  wire ctrl_ready_r;
  wire [4:0] ctrl_opcode_rrrr;
  wire [4:0] ctrl_opcode_rrrrr;
  wire [4:0] ctrl_opcode_rrrrrr;
  wire [4:0] ctrl_opcode_rrrrrrr;
  wire [4:0] ctrl_opcode_rrrrrrrr;
  wire [10:0] ctrl_goto_addr_rrrr;
  wire [10:0] ctrl_goto_addr_rrrrr;
  wire [10:0] ctrl_goto_addr_rrrrrr;
  wire [10:0] ctrl_goto_addr_rrrrrrr;
  wire [10:0] ctrl_goto_addr_rrrrrrrr;
  wire ctrl_jump;
  wire ctrl_ret_func;
  wire [10:0] next_addr;
  wire ready;
  wire [7:0] instruction_pcore_enable_r;
  wire [7:0] instruction_pcore_enable_rr;
  wire tid_vm;
  wire tid_vm_r;
  wire tid_vm_rr;
  wire [1:0] task_data_model;
  wire [1:0] task_data_model_r;
  wire [1:0] task_data_model_rr;
  wire [27:0] tid_iregister_auto;
  wire [27:0] tid_iregister_auto_r;
  wire ready2;
  wire [3:0] n14290_o;
  wire [10:0] n14294_o;
  wire n14296_o;
  wire n14297_o;
  wire n14298_o;
  wire n14299_o;
  wire n14300_o;
  wire n14301_o;
  wire n14304_o;
  wire n14305_o;
  wire n14306_o;
  wire n14307_o;
  wire n14308_o;
  wire n14312_o;
  wire n14313_o;
  wire n14314_o;
  wire n14315_o;
  wire n14316_o;
  wire [15:0] delay_i_n14318;
  localparam n14319_o = 1'b1;
  wire [15:0] delay_i_out_out;
  wire n14325_o;
  wire n14326_o;
  wire n14327_o;
  wire n14328_o;
  wire n14329_o;
  wire n14332_o;
  wire n14333_o;
  wire n14334_o;
  wire n14335_o;
  wire n14336_o;
  wire n14337_o;
  wire n14340_o;
  wire n14341_o;
  wire n14342_o;
  wire n14343_o;
  wire n14344_o;
  wire n14345_o;
  wire n14348_o;
  wire n14349_o;
  wire n14350_o;
  wire n14351_o;
  wire n14352_o;
  wire n14353_o;
  wire n14356_o;
  wire n14357_o;
  wire n14358_o;
  wire n14359_o;
  wire n14360_o;
  wire n14361_o;
  wire n14364_o;
  wire n14365_o;
  wire n14366_o;
  wire n14367_o;
  wire n14368_o;
  wire n14369_o;
  wire n14372_o;
  wire n14373_o;
  wire n14374_o;
  wire n14375_o;
  wire n14376_o;
  wire n14377_o;
  wire n14380_o;
  wire n14381_o;
  wire n14382_o;
  wire n14383_o;
  wire n14384_o;
  wire n14385_o;
  wire n14388_o;
  wire n14389_o;
  wire n14390_o;
  wire n14391_o;
  wire n14392_o;
  wire n14393_o;
  wire n14396_o;
  wire n14397_o;
  wire n14398_o;
  wire n14399_o;
  wire n14400_o;
  wire n14401_o;
  wire n14404_o;
  wire n14405_o;
  wire n14406_o;
  wire n14407_o;
  wire n14408_o;
  wire n14409_o;
  wire n14412_o;
  wire n14413_o;
  wire n14414_o;
  wire n14415_o;
  wire n14416_o;
  wire n14417_o;
  wire n14420_o;
  wire n14421_o;
  wire n14422_o;
  wire n14423_o;
  wire n14424_o;
  wire n14425_o;
  wire n14428_o;
  wire n14429_o;
  wire n14430_o;
  wire n14431_o;
  wire n14432_o;
  wire n14433_o;
  wire n14436_o;
  wire n14437_o;
  wire n14438_o;
  wire n14439_o;
  wire n14440_o;
  wire n14441_o;
  wire n14444_o;
  wire n14445_o;
  wire n14446_o;
  wire n14447_o;
  wire n14448_o;
  wire n14449_o;
  wire n14452_o;
  localparam [1:0] n14453_o = 2'b00;
  wire n14454_o;
  wire n14455_o;
  wire n14456_o;
  wire n14457_o;
  wire n14458_o;
  wire n14459_o;
  localparam [1:0] n14460_o = 2'b00;
  wire n14461_o;
  wire [1:0] n14462_o;
  wire n14463_o;
  wire n14464_o;
  wire n14465_o;
  wire n14466_o;
  wire n14467_o;
  wire [1:0] n14468_o;
  wire n14469_o;
  wire n14470_o;
  wire n14471_o;
  wire n14472_o;
  wire n14473_o;
  wire n14474_o;
  wire [1:0] n14475_o;
  wire n14476_o;
  wire n14477_o;
  wire n14478_o;
  wire n14479_o;
  wire n14480_o;
  wire [1:0] n14481_o;
  wire n14482_o;
  wire n14483_o;
  wire n14484_o;
  wire n14485_o;
  wire n14486_o;
  wire n14487_o;
  wire [1:0] n14488_o;
  wire n14489_o;
  wire n14490_o;
  wire n14491_o;
  wire n14492_o;
  wire n14493_o;
  wire [1:0] n14494_o;
  wire n14495_o;
  wire n14496_o;
  wire n14497_o;
  wire n14498_o;
  wire n14499_o;
  wire n14500_o;
  wire [1:0] n14501_o;
  wire n14502_o;
  wire n14503_o;
  wire n14504_o;
  wire n14505_o;
  wire n14506_o;
  wire [1:0] n14507_o;
  wire n14508_o;
  wire n14509_o;
  wire n14510_o;
  wire n14511_o;
  wire n14512_o;
  wire n14513_o;
  wire [1:0] n14514_o;
  wire n14515_o;
  wire n14516_o;
  wire n14517_o;
  wire n14518_o;
  wire n14519_o;
  wire [1:0] n14520_o;
  wire n14521_o;
  wire n14522_o;
  wire n14523_o;
  wire n14524_o;
  wire n14525_o;
  wire n14526_o;
  wire [1:0] n14527_o;
  wire n14528_o;
  wire n14529_o;
  wire n14530_o;
  wire n14531_o;
  wire n14532_o;
  wire [1:0] n14533_o;
  wire n14534_o;
  wire n14535_o;
  wire n14536_o;
  wire n14537_o;
  wire n14538_o;
  wire n14539_o;
  wire [1:0] n14540_o;
  wire n14541_o;
  wire n14542_o;
  wire n14543_o;
  wire n14544_o;
  wire n14545_o;
  wire [1:0] n14546_o;
  wire n14547_o;
  wire n14548_o;
  wire n14549_o;
  wire n14550_o;
  wire n14551_o;
  wire n14552_o;
  wire [1:0] n14553_o;
  wire n14554_o;
  wire n14555_o;
  wire n14556_o;
  wire n14557_o;
  wire n14558_o;
  wire [1:0] n14559_o;
  wire n14560_o;
  wire n14561_o;
  wire n14562_o;
  wire n14563_o;
  wire n14564_o;
  wire n14565_o;
  wire [1:0] n14566_o;
  wire n14567_o;
  wire n14568_o;
  wire n14569_o;
  wire n14570_o;
  wire n14571_o;
  wire [1:0] n14572_o;
  wire n14573_o;
  wire n14574_o;
  wire n14575_o;
  wire n14576_o;
  wire n14577_o;
  wire n14578_o;
  wire [1:0] n14579_o;
  wire n14580_o;
  wire n14581_o;
  wire n14582_o;
  wire n14583_o;
  wire n14584_o;
  wire [1:0] n14585_o;
  wire n14586_o;
  wire n14587_o;
  wire n14588_o;
  wire n14589_o;
  wire n14590_o;
  wire n14591_o;
  wire [1:0] n14592_o;
  wire n14593_o;
  wire n14594_o;
  wire n14595_o;
  wire n14596_o;
  wire n14597_o;
  wire [1:0] n14598_o;
  wire n14599_o;
  wire n14600_o;
  wire n14601_o;
  wire n14602_o;
  wire n14603_o;
  wire n14604_o;
  wire [1:0] n14605_o;
  wire n14606_o;
  wire n14607_o;
  wire n14608_o;
  wire n14609_o;
  wire n14610_o;
  wire [1:0] n14611_o;
  wire n14612_o;
  wire n14613_o;
  wire n14614_o;
  wire n14615_o;
  wire n14616_o;
  wire n14617_o;
  wire [1:0] n14618_o;
  wire n14619_o;
  wire n14620_o;
  wire n14621_o;
  wire n14622_o;
  wire n14623_o;
  wire [1:0] n14624_o;
  wire n14625_o;
  wire n14626_o;
  wire n14627_o;
  wire n14628_o;
  wire n14629_o;
  wire n14630_o;
  wire [1:0] n14631_o;
  wire n14632_o;
  wire n14633_o;
  wire n14634_o;
  wire n14635_o;
  wire n14636_o;
  wire [1:0] n14637_o;
  wire n14638_o;
  wire n14639_o;
  wire n14640_o;
  wire n14641_o;
  wire n14642_o;
  wire n14643_o;
  wire [1:0] n14644_o;
  wire n14645_o;
  wire n14646_o;
  wire n14647_o;
  wire n14648_o;
  wire n14649_o;
  wire [1:0] n14650_o;
  wire n14651_o;
  wire n14652_o;
  wire n14653_o;
  wire n14654_o;
  wire n14655_o;
  wire n14656_o;
  wire [1:0] n14657_o;
  wire n14658_o;
  wire n14659_o;
  wire n14660_o;
  wire n14661_o;
  wire n14662_o;
  wire [1:0] n14663_o;
  wire n14668_o;
  wire [4:0] n14670_o;
  wire n14672_o;
  wire n14673_o;
  wire n14676_o;
  wire [4:0] n14677_o;
  wire n14679_o;
  wire n14680_o;
  wire n14683_o;
  wire [7:0] n14790_o;
  wire n14792_o;
  wire [3:0] n14793_o;
  wire n14795_o;
  wire n14796_o;
  wire n14797_o;
  wire n14798_o;
  wire [3:0] n14801_o;
  wire [3:0] n14803_o;
  wire [3:0] n14805_o;
  wire n14806_o;
  wire n14807_o;
  wire n14808_o;
  wire [3:0] n14811_o;
  wire [3:0] n14813_o;
  wire [3:0] n14815_o;
  wire [3:0] n14816_o;
  wire [3:0] n14817_o;
  wire n14819_o;
  wire n14820_o;
  wire n14821_o;
  wire n14822_o;
  wire [3:0] n14825_o;
  wire [3:0] n14827_o;
  wire [3:0] n14829_o;
  wire n14830_o;
  wire n14831_o;
  wire n14832_o;
  wire [3:0] n14835_o;
  wire [3:0] n14837_o;
  wire [3:0] n14839_o;
  wire [3:0] n14840_o;
  wire [3:0] n14841_o;
  wire [15:0] arbiter_1_i_n14843;
  wire arbiter_1_i_n14844;
  wire [15:0] arbiter_1_i_gnt_out;
  wire arbiter_1_i_gnt_valid_out;
  wire [15:0] n14849_o;
  wire [15:0] n14850_o;
  wire [15:0] n14851_o;
  wire [15:0] n14852_o;
  wire [15:0] n14853_o;
  wire [15:0] n14854_o;
  wire n14862_o;
  wire n14864_o;
  wire n14866_o;
  wire n14868_o;
  wire n14870_o;
  wire n14872_o;
  wire n14874_o;
  wire n14876_o;
  wire n14878_o;
  wire n14880_o;
  wire n14882_o;
  wire n14884_o;
  wire n14886_o;
  wire n14888_o;
  wire n14890_o;
  wire [14:0] n14891_o;
  reg [15:0] n14908_o;
  wire n14918_o;
  wire [4:0] n14923_o;
  wire n14931_o;
  wire n14932_o;
  wire n14933_o;
  wire n14934_o;
  wire n14935_o;
  wire n14937_o;
  wire n14938_o;
  wire [4:0] n14940_o;
  wire [4:0] n14941_o;
  wire n14943_o;
  wire n14944_o;
  wire n14945_o;
  wire n14946_o;
  wire n14947_o;
  wire n14948_o;
  wire n14949_o;
  wire n14951_o;
  wire n14952_o;
  wire n14953_o;
  wire n14955_o;
  wire n14957_o;
  wire n14958_o;
  wire [1:0] n14959_o;
  wire n14960_o;
  wire n14961_o;
  wire [10:0] n14962_o;
  wire n14963_o;
  wire n14964_o;
  wire n14965_o;
  wire n14966_o;
  wire n14968_o;
  wire n14970_o;
  wire [10:0] n14971_o;
  wire n14972_o;
  wire n14974_o;
  wire n14975_o;
  wire n14976_o;
  wire n14977_o;
  wire n14978_o;
  wire n14979_o;
  wire n14980_o;
  wire [10:0] n14986_o;
  wire n14988_o;
  wire n14989_o;
  wire n14990_o;
  wire [1:0] n14991_o;
  wire n14994_o;
  wire [27:0] n14995_o;
  wire [27:0] n14996_o;
  wire n14997_o;
  wire n14998_o;
  wire n14999_o;
  wire n15000_o;
  wire n15001_o;
  wire n15004_o;
  wire n15005_o;
  wire n15006_o;
  wire n15007_o;
  wire n15008_o;
  wire n15009_o;
  wire n15010_o;
  wire n15011_o;
  wire n15013_o;
  wire n15014_o;
  wire n15015_o;
  wire n15017_o;
  wire n15019_o;
  wire n15020_o;
  wire [1:0] n15021_o;
  wire n15022_o;
  wire n15023_o;
  wire [10:0] n15024_o;
  wire n15025_o;
  wire n15026_o;
  wire n15027_o;
  wire n15028_o;
  wire n15030_o;
  wire n15032_o;
  wire [10:0] n15033_o;
  wire n15034_o;
  wire n15036_o;
  wire n15037_o;
  wire n15038_o;
  wire n15039_o;
  wire n15040_o;
  wire n15041_o;
  wire n15042_o;
  wire [10:0] n15048_o;
  wire n15050_o;
  wire n15051_o;
  wire n15052_o;
  wire [1:0] n15053_o;
  wire n15056_o;
  wire [27:0] n15057_o;
  wire [27:0] n15058_o;
  wire n15059_o;
  wire n15060_o;
  wire n15061_o;
  wire n15062_o;
  wire n15063_o;
  wire n15066_o;
  wire n15067_o;
  wire n15068_o;
  wire n15069_o;
  wire n15070_o;
  wire n15071_o;
  wire n15072_o;
  wire n15073_o;
  wire n15075_o;
  wire n15076_o;
  wire n15077_o;
  wire n15079_o;
  wire n15081_o;
  wire n15082_o;
  wire [1:0] n15083_o;
  wire n15084_o;
  wire n15085_o;
  wire [10:0] n15086_o;
  wire n15087_o;
  wire n15088_o;
  wire n15089_o;
  wire n15090_o;
  wire n15092_o;
  wire n15094_o;
  wire [10:0] n15095_o;
  wire n15096_o;
  wire n15098_o;
  wire n15099_o;
  wire n15100_o;
  wire n15101_o;
  wire n15102_o;
  wire n15103_o;
  wire n15104_o;
  wire [10:0] n15110_o;
  wire n15112_o;
  wire n15113_o;
  wire n15114_o;
  wire [1:0] n15115_o;
  wire n15118_o;
  wire [27:0] n15119_o;
  wire [27:0] n15120_o;
  wire n15121_o;
  wire n15122_o;
  wire n15123_o;
  wire n15124_o;
  wire n15125_o;
  wire n15128_o;
  wire n15129_o;
  wire n15130_o;
  wire n15131_o;
  wire n15132_o;
  wire n15133_o;
  wire n15134_o;
  wire n15135_o;
  wire n15137_o;
  wire n15138_o;
  wire n15139_o;
  wire n15141_o;
  wire n15143_o;
  wire n15144_o;
  wire [1:0] n15145_o;
  wire n15146_o;
  wire n15147_o;
  wire [10:0] n15148_o;
  wire n15149_o;
  wire n15150_o;
  wire n15151_o;
  wire n15152_o;
  wire n15154_o;
  wire n15156_o;
  wire [10:0] n15157_o;
  wire n15158_o;
  wire n15160_o;
  wire n15161_o;
  wire n15162_o;
  wire n15163_o;
  wire n15164_o;
  wire n15165_o;
  wire n15166_o;
  wire [10:0] n15172_o;
  wire n15174_o;
  wire n15175_o;
  wire n15176_o;
  wire [1:0] n15177_o;
  wire n15180_o;
  wire [27:0] n15181_o;
  wire [27:0] n15182_o;
  wire n15183_o;
  wire n15184_o;
  wire n15185_o;
  wire n15186_o;
  wire n15187_o;
  wire n15190_o;
  wire n15191_o;
  wire n15192_o;
  wire n15193_o;
  wire n15194_o;
  wire n15195_o;
  wire n15196_o;
  wire n15197_o;
  wire n15199_o;
  wire n15200_o;
  wire n15201_o;
  wire n15203_o;
  wire n15205_o;
  wire n15206_o;
  wire [1:0] n15207_o;
  wire n15208_o;
  wire n15209_o;
  wire [10:0] n15210_o;
  wire n15211_o;
  wire n15212_o;
  wire n15213_o;
  wire n15214_o;
  wire n15216_o;
  wire n15218_o;
  wire [10:0] n15219_o;
  wire n15220_o;
  wire n15222_o;
  wire n15223_o;
  wire n15224_o;
  wire n15225_o;
  wire n15226_o;
  wire n15227_o;
  wire n15228_o;
  wire [10:0] n15234_o;
  wire n15236_o;
  wire n15237_o;
  wire n15238_o;
  wire [1:0] n15239_o;
  wire n15242_o;
  wire [27:0] n15243_o;
  wire [27:0] n15244_o;
  wire n15245_o;
  wire n15246_o;
  wire n15247_o;
  wire n15248_o;
  wire n15249_o;
  wire n15252_o;
  wire n15253_o;
  wire n15254_o;
  wire n15255_o;
  wire n15256_o;
  wire n15257_o;
  wire n15258_o;
  wire n15259_o;
  wire n15261_o;
  wire n15262_o;
  wire n15263_o;
  wire n15265_o;
  wire n15267_o;
  wire n15268_o;
  wire [1:0] n15269_o;
  wire n15270_o;
  wire n15271_o;
  wire [10:0] n15272_o;
  wire n15273_o;
  wire n15274_o;
  wire n15275_o;
  wire n15276_o;
  wire n15278_o;
  wire n15280_o;
  wire [10:0] n15281_o;
  wire n15282_o;
  wire n15284_o;
  wire n15285_o;
  wire n15286_o;
  wire n15287_o;
  wire n15288_o;
  wire n15289_o;
  wire n15290_o;
  wire [10:0] n15296_o;
  wire n15298_o;
  wire n15299_o;
  wire n15300_o;
  wire [1:0] n15301_o;
  wire n15304_o;
  wire [27:0] n15305_o;
  wire [27:0] n15306_o;
  wire n15307_o;
  wire n15308_o;
  wire n15309_o;
  wire n15310_o;
  wire n15311_o;
  wire n15314_o;
  wire n15315_o;
  wire n15316_o;
  wire n15317_o;
  wire n15318_o;
  wire n15319_o;
  wire n15320_o;
  wire n15321_o;
  wire n15323_o;
  wire n15324_o;
  wire n15325_o;
  wire n15327_o;
  wire n15329_o;
  wire n15330_o;
  wire [1:0] n15331_o;
  wire n15332_o;
  wire n15333_o;
  wire [10:0] n15334_o;
  wire n15335_o;
  wire n15336_o;
  wire n15337_o;
  wire n15338_o;
  wire n15340_o;
  wire n15342_o;
  wire [10:0] n15343_o;
  wire n15344_o;
  wire n15346_o;
  wire n15347_o;
  wire n15348_o;
  wire n15349_o;
  wire n15350_o;
  wire n15351_o;
  wire n15352_o;
  wire [10:0] n15358_o;
  wire n15360_o;
  wire n15361_o;
  wire n15362_o;
  wire [1:0] n15363_o;
  wire n15366_o;
  wire [27:0] n15367_o;
  wire [27:0] n15368_o;
  wire n15369_o;
  wire n15370_o;
  wire n15371_o;
  wire n15372_o;
  wire n15373_o;
  wire n15376_o;
  wire n15377_o;
  wire n15378_o;
  wire n15379_o;
  wire n15380_o;
  wire n15381_o;
  wire n15382_o;
  wire n15383_o;
  wire n15385_o;
  wire n15386_o;
  wire n15387_o;
  wire n15389_o;
  wire n15391_o;
  wire n15392_o;
  wire [1:0] n15393_o;
  wire n15394_o;
  wire n15395_o;
  wire [10:0] n15396_o;
  wire n15397_o;
  wire n15398_o;
  wire n15399_o;
  wire n15400_o;
  wire n15402_o;
  wire n15404_o;
  wire [10:0] n15405_o;
  wire n15406_o;
  wire n15408_o;
  wire n15409_o;
  wire n15410_o;
  wire n15411_o;
  wire n15412_o;
  wire n15413_o;
  wire n15414_o;
  wire [10:0] n15420_o;
  wire n15422_o;
  wire n15423_o;
  wire n15424_o;
  wire [1:0] n15425_o;
  wire n15428_o;
  wire [27:0] n15429_o;
  wire [27:0] n15430_o;
  wire n15431_o;
  wire n15432_o;
  wire n15433_o;
  wire n15434_o;
  wire n15435_o;
  wire n15438_o;
  wire n15439_o;
  wire n15440_o;
  wire n15441_o;
  wire n15442_o;
  wire n15443_o;
  wire n15444_o;
  wire n15445_o;
  wire n15447_o;
  wire n15448_o;
  wire n15449_o;
  wire n15451_o;
  wire n15453_o;
  wire n15454_o;
  wire [1:0] n15455_o;
  wire n15456_o;
  wire n15457_o;
  wire [10:0] n15458_o;
  wire n15459_o;
  wire n15460_o;
  wire n15461_o;
  wire n15462_o;
  wire n15464_o;
  wire n15466_o;
  wire [10:0] n15467_o;
  wire n15468_o;
  wire n15470_o;
  wire n15471_o;
  wire n15472_o;
  wire n15473_o;
  wire n15474_o;
  wire n15475_o;
  wire n15476_o;
  wire [10:0] n15482_o;
  wire n15484_o;
  wire n15485_o;
  wire n15486_o;
  wire [1:0] n15487_o;
  wire n15490_o;
  wire [27:0] n15491_o;
  wire [27:0] n15492_o;
  wire n15493_o;
  wire n15494_o;
  wire n15495_o;
  wire n15496_o;
  wire n15497_o;
  wire n15500_o;
  wire n15501_o;
  wire n15502_o;
  wire n15503_o;
  wire n15504_o;
  wire n15505_o;
  wire n15506_o;
  wire n15507_o;
  wire n15509_o;
  wire n15510_o;
  wire n15511_o;
  wire n15513_o;
  wire n15515_o;
  wire n15516_o;
  wire [1:0] n15517_o;
  wire n15518_o;
  wire n15519_o;
  wire [10:0] n15520_o;
  wire n15521_o;
  wire n15522_o;
  wire n15523_o;
  wire n15524_o;
  wire n15526_o;
  wire n15528_o;
  wire [10:0] n15529_o;
  wire n15530_o;
  wire n15532_o;
  wire n15533_o;
  wire n15534_o;
  wire n15535_o;
  wire n15536_o;
  wire n15537_o;
  wire n15538_o;
  wire [10:0] n15544_o;
  wire n15546_o;
  wire n15547_o;
  wire n15548_o;
  wire [1:0] n15549_o;
  wire n15552_o;
  wire [27:0] n15553_o;
  wire [27:0] n15554_o;
  wire n15555_o;
  wire n15556_o;
  wire n15557_o;
  wire n15558_o;
  wire n15559_o;
  wire n15562_o;
  wire n15563_o;
  wire n15564_o;
  wire n15565_o;
  wire n15566_o;
  wire n15567_o;
  wire n15568_o;
  wire n15569_o;
  wire n15571_o;
  wire n15572_o;
  wire n15573_o;
  wire n15575_o;
  wire n15577_o;
  wire n15578_o;
  wire [1:0] n15579_o;
  wire n15580_o;
  wire n15581_o;
  wire [10:0] n15582_o;
  wire n15583_o;
  wire n15584_o;
  wire n15585_o;
  wire n15586_o;
  wire n15588_o;
  wire n15590_o;
  wire [10:0] n15591_o;
  wire n15592_o;
  wire n15594_o;
  wire n15595_o;
  wire n15596_o;
  wire n15597_o;
  wire n15598_o;
  wire n15599_o;
  wire n15600_o;
  wire [10:0] n15606_o;
  wire n15608_o;
  wire n15609_o;
  wire n15610_o;
  wire [1:0] n15611_o;
  wire n15614_o;
  wire [27:0] n15615_o;
  wire [27:0] n15616_o;
  wire n15617_o;
  wire n15618_o;
  wire n15619_o;
  wire n15620_o;
  wire n15621_o;
  wire n15624_o;
  wire n15625_o;
  wire n15626_o;
  wire n15627_o;
  wire n15628_o;
  wire n15629_o;
  wire n15630_o;
  wire n15631_o;
  wire n15633_o;
  wire n15634_o;
  wire n15635_o;
  wire n15637_o;
  wire n15639_o;
  wire n15640_o;
  wire [1:0] n15641_o;
  wire n15642_o;
  wire n15643_o;
  wire [10:0] n15644_o;
  wire n15645_o;
  wire n15646_o;
  wire n15647_o;
  wire n15648_o;
  wire n15650_o;
  wire n15652_o;
  wire [10:0] n15653_o;
  wire n15654_o;
  wire n15656_o;
  wire n15657_o;
  wire n15658_o;
  wire n15659_o;
  wire n15660_o;
  wire n15661_o;
  wire n15662_o;
  wire [10:0] n15668_o;
  wire n15670_o;
  wire n15671_o;
  wire n15672_o;
  wire [1:0] n15673_o;
  wire n15676_o;
  wire [27:0] n15677_o;
  wire [27:0] n15678_o;
  wire n15679_o;
  wire n15680_o;
  wire n15681_o;
  wire n15682_o;
  wire n15683_o;
  wire n15686_o;
  wire n15687_o;
  wire n15688_o;
  wire n15689_o;
  wire n15690_o;
  wire n15691_o;
  wire n15692_o;
  wire n15693_o;
  wire n15695_o;
  wire n15696_o;
  wire n15697_o;
  wire n15699_o;
  wire n15701_o;
  wire n15702_o;
  wire [1:0] n15703_o;
  wire n15704_o;
  wire n15705_o;
  wire [10:0] n15706_o;
  wire n15707_o;
  wire n15708_o;
  wire n15709_o;
  wire n15710_o;
  wire n15712_o;
  wire n15714_o;
  wire [10:0] n15715_o;
  wire n15716_o;
  wire n15718_o;
  wire n15719_o;
  wire n15720_o;
  wire n15721_o;
  wire n15722_o;
  wire n15723_o;
  wire n15724_o;
  wire [10:0] n15730_o;
  wire n15732_o;
  wire n15733_o;
  wire n15734_o;
  wire [1:0] n15735_o;
  wire n15738_o;
  wire [27:0] n15739_o;
  wire [27:0] n15740_o;
  wire n15741_o;
  wire n15742_o;
  wire n15743_o;
  wire n15744_o;
  wire n15745_o;
  wire n15748_o;
  wire n15749_o;
  wire n15750_o;
  wire n15751_o;
  wire n15752_o;
  wire n15753_o;
  wire n15754_o;
  wire n15755_o;
  wire n15757_o;
  wire n15758_o;
  wire n15759_o;
  wire n15761_o;
  wire n15763_o;
  wire n15764_o;
  wire [1:0] n15765_o;
  wire n15766_o;
  wire n15767_o;
  wire [10:0] n15768_o;
  wire n15769_o;
  wire n15770_o;
  wire n15771_o;
  wire n15772_o;
  wire n15774_o;
  wire n15776_o;
  wire [10:0] n15777_o;
  wire n15778_o;
  wire n15780_o;
  wire n15781_o;
  wire n15782_o;
  wire n15783_o;
  wire n15784_o;
  wire n15785_o;
  wire n15786_o;
  wire [10:0] n15792_o;
  wire n15794_o;
  wire n15795_o;
  wire n15796_o;
  wire [1:0] n15797_o;
  wire n15800_o;
  wire [27:0] n15801_o;
  wire [27:0] n15802_o;
  wire n15803_o;
  wire n15804_o;
  wire n15805_o;
  wire n15806_o;
  wire n15807_o;
  wire n15810_o;
  wire n15811_o;
  wire n15812_o;
  wire n15813_o;
  wire n15814_o;
  wire n15815_o;
  wire n15816_o;
  wire n15817_o;
  wire n15819_o;
  wire n15820_o;
  wire n15821_o;
  wire n15823_o;
  wire n15825_o;
  wire n15826_o;
  wire [1:0] n15827_o;
  wire n15828_o;
  wire n15829_o;
  wire [10:0] n15830_o;
  wire n15831_o;
  wire n15832_o;
  wire n15833_o;
  wire n15834_o;
  wire n15836_o;
  wire n15838_o;
  wire [10:0] n15839_o;
  wire n15840_o;
  wire n15842_o;
  wire n15843_o;
  wire n15844_o;
  wire n15845_o;
  wire n15846_o;
  wire n15847_o;
  wire n15848_o;
  wire n15849_o;
  wire n15850_o;
  wire n15851_o;
  wire n15852_o;
  wire n15853_o;
  wire [10:0] n15854_o;
  wire n15856_o;
  wire n15857_o;
  wire n15858_o;
  wire [1:0] n15859_o;
  wire n15862_o;
  wire [27:0] n15863_o;
  wire [27:0] n15864_o;
  wire n15865_o;
  wire n15866_o;
  wire n15867_o;
  wire n15868_o;
  wire n15869_o;
  wire n15872_o;
  wire n15873_o;
  wire n15874_o;
  wire n15875_o;
  wire n15876_o;
  wire n15877_o;
  wire n15878_o;
  wire n15879_o;
  wire n15881_o;
  wire n15882_o;
  wire n15883_o;
  wire n15885_o;
  wire n15887_o;
  wire n15888_o;
  wire [1:0] n15889_o;
  wire n15890_o;
  wire n15891_o;
  wire [10:0] n15892_o;
  wire n15893_o;
  wire n15894_o;
  wire n15895_o;
  wire n15896_o;
  wire n15898_o;
  wire n15900_o;
  wire [10:0] n15901_o;
  wire n15902_o;
  wire n15904_o;
  wire n15905_o;
  wire [10:0] n15906_o;
  wire n15908_o;
  wire n15909_o;
  wire n15910_o;
  wire [1:0] n15911_o;
  wire n15914_o;
  wire [27:0] n15915_o;
  wire [27:0] n15916_o;
  wire n15917_o;
  wire n15918_o;
  wire n15919_o;
  wire n15920_o;
  wire n15921_o;
  wire n15924_o;
  wire [175:0] n15925_o;
  wire [15:0] n15927_o;
  wire [15:0] n15929_o;
  wire [31:0] n15932_o;
  wire [447:0] n15935_o;
  wire [15:0] n15938_o;
  wire [15:0] n15940_o;
  wire [15:0] n15947_o;
  wire [79:0] n16036_o;
  wire [31:0] n16037_o;
  wire [15:0] n16038_o;
  wire n16042_o;
  wire [4:0] n16044_o;
  wire n16046_o;
  wire n16047_o;
  wire n16050_o;
  wire [4:0] n16051_o;
  wire [10:0] n16052_o;
  wire [9:0] n16053_o;
  wire [9:0] n16055_o;
  wire [10:0] n16057_o;
  wire [10:0] n16059_o;
  wire n16061_o;
  wire n16062_o;
  wire n16065_o;
  wire [10:0] n16080_o;
  wire n16161_o;
  wire n16163_o;
  wire n16164_o;
  wire n16166_o;
  wire n16167_o;
  wire n16168_o;
  wire n16169_o;
  wire n16171_o;
  wire n16172_o;
  wire n16174_o;
  wire n16176_o;
  wire n16177_o;
  wire n16179_o;
  wire n16181_o;
  wire [7:0] n16182_o;
  reg n16186_o;
  reg n16196_o;
  wire n16198_o;
  wire n16200_o;
  wire n16204_o;
  wire n16215_o;
  wire n16217_o;
  wire n16219_o;
  wire n16222_o;
  wire n16224_o;
  wire n16227_o;
  wire n16229_o;
  wire n16232_o;
  wire n16234_o;
  wire n16237_o;
  wire n16239_o;
  wire n16242_o;
  wire n16244_o;
  wire n16247_o;
  wire n16249_o;
  wire n16252_o;
  wire n16254_o;
  wire n16257_o;
  wire n16259_o;
  wire n16262_o;
  wire n16264_o;
  wire n16267_o;
  wire n16269_o;
  wire n16272_o;
  wire n16274_o;
  wire n16277_o;
  wire n16279_o;
  wire n16282_o;
  wire n16284_o;
  wire n16287_o;
  wire n16289_o;
  wire n16292_o;
  wire n16294_o;
  wire n16297_o;
  wire [7:0] n16298_o;
  wire [7:0] n16299_o;
  wire [7:0] n16300_o;
  reg [175:0] n16308_q;
  reg [15:0] n16309_q;
  reg [15:0] n16310_q;
  reg [15:0] n16311_q;
  reg [31:0] n16312_q;
  reg [31:0] n16313_q;
  reg [447:0] n16314_q;
  reg [447:0] n16315_q;
  reg [15:0] n16325_q;
  reg n16326_q;
  reg [15:0] n16327_q;
  reg n16328_q;
  reg n16329_q;
  reg [15:0] n16330_q;
  reg [15:0] n16331_q;
  reg [15:0] n16332_q;
  reg [15:0] n16333_q;
  reg [15:0] n16334_q;
  reg [15:0] n16335_q;
  reg [15:0] n16336_q;
  reg [15:0] n16337_q;
  reg [15:0] n16338_q;
  reg [3:0] n16339_q;
  reg [3:0] n16340_q;
  reg [3:0] n16341_q;
  reg [10:0] n16342_q;
  reg [10:0] n16343_q;
  reg [15:0] n16344_q;
  wire [15:0] n16345_o;
  reg [1:0] n16346_q;
  reg [15:0] n16347_q;
  reg [79:0] n16348_q;
  reg [31:0] n16349_q;
  reg n16350_q;
  reg n16351_q;
  wire [10:0] n16352_o;
  reg [10:0] n16353_q;
  wire [4:0] n16354_o;
  reg [4:0] n16355_q;
  reg [4:0] n16356_q;
  wire [15:0] n16357_o;
  reg [15:0] n16358_q;
  wire n16359_o;
  reg n16360_q;
  reg [15:0] n16361_q;
  wire n16362_o;
  reg n16363_q;
  wire [27:0] n16364_o;
  reg [27:0] n16365_q;
  wire [1:0] n16366_o;
  reg [1:0] n16367_q;
  reg [10:0] n16368_q;
  reg [10:0] n16369_q;
  wire n16370_o;
  wire n16371_o;
  reg n16372_q;
  reg n16373_q;
  reg n16374_q;
  reg n16375_q;
  reg n16376_q;
  reg n16377_q;
  reg n16378_q;
  reg n16379_q;
  wire n16380_o;
  wire [4:0] n16381_o;
  reg [4:0] n16382_q;
  wire n16383_o;
  wire [10:0] n16384_o;
  reg [10:0] n16385_q;
  reg [4:0] n16386_q;
  reg [10:0] n16387_q;
  reg [4:0] n16388_q;
  reg [10:0] n16389_q;
  reg [10:0] n16390_q;
  reg [10:0] n16391_q;
  reg [10:0] n16392_q;
  reg [10:0] n16393_q;
  reg [10:0] n16394_q;
  reg [10:0] n16395_q;
  reg n16396_q;
  reg [4:0] n16397_q;
  reg [4:0] n16398_q;
  reg [4:0] n16399_q;
  reg [4:0] n16400_q;
  reg [4:0] n16401_q;
  reg [10:0] n16402_q;
  reg [10:0] n16403_q;
  reg [10:0] n16404_q;
  reg [10:0] n16405_q;
  reg [10:0] n16406_q;
  reg [7:0] n16407_q;
  reg [7:0] n16408_q;
  reg n16409_q;
  reg n16410_q;
  reg [1:0] n16411_q;
  reg [1:0] n16412_q;
  reg [27:0] n16413_q;
  wire [1:0] n16414_o;
  wire [27:0] n16415_o;
  wire [27:0] n16416_o;
  wire [27:0] n16417_o;
  wire [27:0] n16418_o;
  wire [27:0] n16419_o;
  wire [27:0] n16420_o;
  wire [27:0] n16421_o;
  wire [27:0] n16422_o;
  wire [27:0] n16423_o;
  wire [27:0] n16424_o;
  wire [27:0] n16425_o;
  wire [27:0] n16426_o;
  wire [27:0] n16427_o;
  wire [27:0] n16428_o;
  wire [27:0] n16429_o;
  wire [27:0] n16430_o;
  wire [1:0] n16431_o;
  reg [27:0] n16432_o;
  wire [1:0] n16433_o;
  reg [27:0] n16434_o;
  wire [1:0] n16435_o;
  reg [27:0] n16436_o;
  wire [1:0] n16437_o;
  reg [27:0] n16438_o;
  wire [1:0] n16439_o;
  reg [27:0] n16440_o;
  wire n16441_o;
  wire n16442_o;
  wire n16443_o;
  wire n16444_o;
  wire n16445_o;
  wire n16446_o;
  wire n16447_o;
  wire n16448_o;
  wire n16449_o;
  wire n16450_o;
  wire n16451_o;
  wire n16452_o;
  wire n16453_o;
  wire n16454_o;
  wire n16455_o;
  wire n16456_o;
  wire [1:0] n16457_o;
  reg n16458_o;
  wire [1:0] n16459_o;
  reg n16460_o;
  wire [1:0] n16461_o;
  reg n16462_o;
  wire [1:0] n16463_o;
  reg n16464_o;
  wire [1:0] n16465_o;
  reg n16466_o;
  wire [1:0] n16467_o;
  wire [1:0] n16468_o;
  wire [1:0] n16469_o;
  wire [1:0] n16470_o;
  wire [1:0] n16471_o;
  wire [1:0] n16472_o;
  wire [1:0] n16473_o;
  wire [1:0] n16474_o;
  wire [1:0] n16475_o;
  wire [1:0] n16476_o;
  wire [1:0] n16477_o;
  wire [1:0] n16478_o;
  wire [1:0] n16479_o;
  wire [1:0] n16480_o;
  wire [1:0] n16481_o;
  wire [1:0] n16482_o;
  wire [1:0] n16483_o;
  reg [1:0] n16484_o;
  wire [1:0] n16485_o;
  reg [1:0] n16486_o;
  wire [1:0] n16487_o;
  reg [1:0] n16488_o;
  wire [1:0] n16489_o;
  reg [1:0] n16490_o;
  wire [1:0] n16491_o;
  reg [1:0] n16492_o;
  wire [10:0] n16493_o;
  wire [10:0] n16494_o;
  wire [10:0] n16495_o;
  wire [10:0] n16496_o;
  wire [10:0] n16497_o;
  wire [10:0] n16498_o;
  wire [10:0] n16499_o;
  wire [10:0] n16500_o;
  wire [10:0] n16501_o;
  wire [10:0] n16502_o;
  wire [10:0] n16503_o;
  wire [10:0] n16504_o;
  wire [10:0] n16505_o;
  wire [10:0] n16506_o;
  wire [10:0] n16507_o;
  wire [10:0] n16508_o;
  wire [1:0] n16509_o;
  reg [10:0] n16510_o;
  wire [1:0] n16511_o;
  reg [10:0] n16512_o;
  wire [1:0] n16513_o;
  reg [10:0] n16514_o;
  wire [1:0] n16515_o;
  reg [10:0] n16516_o;
  wire [1:0] n16517_o;
  reg [10:0] n16518_o;
  assign instruction_mu_out = instruction_mu_r;
  assign instruction_imu_out = instruction_imu_r;
  assign instruction_mu_valid_out = instruction_mu_valid_r;
  assign instruction_imu_valid_out = instruction_imu_valid_r;
  assign instruction_vm_out = tid_vm_rr;
  assign instruction_data_model_out = task_data_model_rr;
  assign instruction_tid_out = tid2_rrr;
  assign instruction_tid_valid_out = tid_valid_rrr;
  assign instruction_pre_tid_out = tid2_rr;
  assign instruction_pre_tid_valid_out = tid_valid_rr;
  assign instruction_pre_pre_tid_out = tid2_r;
  assign instruction_pre_pre_tid_valid_out = tid_valid_r;
  assign instruction_pre_pre_vm_out = tid_vm;
  assign instruction_pre_pre_data_model_out = task_data_model;
  assign instruction_pcore_enable_out = instruction_pcore_enable_rr;
  assign instruction_pre_iregister_auto_out = tid_iregister_auto_r;
  assign rom_addr_out = rom_addr;
  assign rom_addr_plus_2_out = n14294_o;
  assign busy_out = n16414_o;
  assign ready_out = ready2;
  /* ../../HW/src/pcore/instr_fetch.vhd:92:8  */
  assign pc_r = n16308_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:93:8  */
  assign busy_r = n16309_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:94:8  */
  assign vm_r = n16310_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:95:8  */
  assign vm_rr = n16311_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:96:8  */
  assign data_model_r = n16312_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:97:8  */
  assign data_model_rr = n16313_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:98:8  */
  assign iregister_auto_r = n16314_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:99:8  */
  assign iregister_auto_rr = n16315_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:109:8  */
  assign tid = n14854_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:110:8  */
  assign tid_delay = delay_i_n14318; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:111:8  */
  assign tid_r = n16325_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:112:8  */
  assign tid_valid_r = n16326_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:113:8  */
  assign tid_rr = n16327_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:114:8  */
  assign tid_valid_rr = n16328_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:115:8  */
  assign tid_valid_rrr = n16329_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:116:8  */
  assign tid_rrr = n16330_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:117:8  */
  assign tid_rrrr = n16331_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:118:8  */
  assign tid_rrrrr = n16332_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:119:8  */
  assign tid_rrrrrr = n16333_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:120:8  */
  assign tid_rrrrrrr = n16334_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:121:8  */
  assign tid_rrrrrrrr = n16335_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:122:8  */
  assign tid_rrrrrrrrr = n16336_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:123:8  */
  assign tid_rrrrrrrrrr = n16337_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:124:8  */
  assign tid_rrrrrrrrrrr = n16338_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:125:8  */
  assign tid2_r = n16339_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:126:8  */
  assign tid2_rr = n16340_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:127:8  */
  assign tid2_rrr = n16341_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:131:8  */
  assign rom_addr = n16518_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:132:8  */
  assign rom_addr_r = n16342_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:133:8  */
  assign rom_addr_rr = n16343_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:138:8  */
  assign delay_r = n16344_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:141:8  */
  assign busy1 = n16345_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:142:8  */
  assign busy2 = n14663_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:143:8  */
  assign busy2_r = n16346_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:147:8  */
  assign avail = avail_r; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:148:8  */
  assign avail_r = n16347_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:149:8  */
  assign next_tid = arbiter_1_i_n14843; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:150:8  */
  assign next_tid2 = n14841_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:151:8  */
  assign next_tid_valid = arbiter_1_i_n14844; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:153:8  */
  assign instruction_mu_r = n16348_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:154:8  */
  assign instruction_imu_r = n16349_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:155:8  */
  assign instruction_mu_valid_r = n16350_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:156:8  */
  assign instruction_imu_valid_r = n16351_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:164:8  */
  assign task_start_addr_r = n16353_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:165:8  */
  assign task_pcore_max_r = n16355_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:166:8  */
  assign task_pcore_curr_r = n16356_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:167:8  */
  always @*
    task_tid_mask_r = n16358_q; // (isignal)
  initial
    task_tid_mask_r = 16'b1111111111111111;
  /* ../../HW/src/pcore/instr_fetch.vhd:168:8  */
  assign task_tid_mask = n14908_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:169:8  */
  assign task_lockstep_r = n16360_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:170:8  */
  assign task_mask_r = n16361_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:171:8  */
  assign task_vm_r = n16363_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:172:8  */
  assign task_iregister_auto_r = n16365_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:173:8  */
  assign task2_data_model_r = n16367_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:175:8  */
  assign mu_instruction = n16036_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:176:8  */
  assign imu_instruction = n16037_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:177:8  */
  assign ctrl_instruction = n16038_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:183:8  */
  assign instruction_addr_r = n16368_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:184:8  */
  assign instruction_addr_rr = n16369_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:186:8  */
  assign got_control_r = n16372_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:187:8  */
  assign got_control_rr = n16373_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:188:8  */
  assign got_control_rrr = n16374_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:189:8  */
  assign got_control_rrrr = n16375_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:190:8  */
  assign got_control_rrrrr = n16376_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:191:8  */
  assign got_control_rrrrrr = n16377_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:192:8  */
  assign got_control_rrrrrrr = n16378_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:193:8  */
  assign got_control_rrrrrrrr = n16379_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:195:8  */
  assign ctrl_opcode_r = n16382_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:196:8  */
  assign ctrl_goto_addr_r = n16385_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:197:8  */
  assign ctrl_opcode_rr = n16386_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:198:8  */
  assign ctrl_goto_addr_rr = n16387_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:199:8  */
  assign ctrl_opcode_rrr = n16388_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:200:8  */
  assign ctrl_goto_addr_rrr = n16389_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:201:8  */
  assign ctrl_next_addr_r = n16390_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:202:8  */
  assign ctrl_next_addr_rr = n16391_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:203:8  */
  assign ctrl_next_addr_rrr = n16392_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:204:8  */
  assign ctrl_next_addr_rrrr = n16393_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:205:8  */
  assign ctrl_next_addr_rrrrr = n16394_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:206:8  */
  assign ctrl_next_addr_rrrrrr = n16395_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:207:8  */
  assign ctrl_ready_r = n16396_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:208:8  */
  assign ctrl_opcode_rrrr = n16397_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:209:8  */
  assign ctrl_opcode_rrrrr = n16398_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:210:8  */
  assign ctrl_opcode_rrrrrr = n16399_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:211:8  */
  assign ctrl_opcode_rrrrrrr = n16400_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:212:8  */
  assign ctrl_opcode_rrrrrrrr = n16401_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:214:8  */
  assign ctrl_goto_addr_rrrr = n16402_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:215:8  */
  assign ctrl_goto_addr_rrrrr = n16403_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:216:8  */
  assign ctrl_goto_addr_rrrrrr = n16404_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:217:8  */
  assign ctrl_goto_addr_rrrrrrr = n16405_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:218:8  */
  assign ctrl_goto_addr_rrrrrrrr = n16406_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:220:8  */
  assign ctrl_jump = n16198_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:221:8  */
  assign ctrl_ret_func = n16200_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:223:8  */
  assign next_addr = ctrl_next_addr_rrrrrr; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:224:8  */
  assign ready = ctrl_ready_r; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:226:8  */
  assign instruction_pcore_enable_r = n16407_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:227:8  */
  assign instruction_pcore_enable_rr = n16408_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:229:8  */
  assign tid_vm = n16466_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:230:8  */
  assign tid_vm_r = n16409_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:231:8  */
  assign tid_vm_rr = n16410_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:233:8  */
  assign task_data_model = n16492_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:234:8  */
  assign task_data_model_r = n16411_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:235:8  */
  assign task_data_model_rr = n16412_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:237:8  */
  assign tid_iregister_auto = n16440_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:238:8  */
  assign tid_iregister_auto_r = n16413_q; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:240:8  */
  assign ready2 = n14316_o; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:366:18  */
  assign n14290_o = 4'b1111 - tid2_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:370:59  */
  assign n14294_o = rom_addr + 11'b00000000010;
  /* ../../HW/src/pcore/instr_fetch.vhd:372:32  */
  assign n14296_o = busy2_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:372:50  */
  assign n14297_o = ~ready2;
  /* ../../HW/src/pcore/instr_fetch.vhd:372:68  */
  assign n14298_o = ~task_vm_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:372:55  */
  assign n14299_o = n14298_o & n14297_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:372:40  */
  assign n14300_o = n14296_o | n14299_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:372:20  */
  assign n14301_o = n14300_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:374:32  */
  assign n14304_o = busy2_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:374:50  */
  assign n14305_o = ~ready2;
  /* ../../HW/src/pcore/instr_fetch.vhd:374:55  */
  assign n14306_o = task_vm_r & n14305_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:374:40  */
  assign n14307_o = n14304_o | n14306_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:374:20  */
  assign n14308_o = n14307_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:376:32  */
  assign n14312_o = task_mask_r == 16'b0000000000000000;
  /* ../../HW/src/pcore/instr_fetch.vhd:377:41  */
  assign n14313_o = task_pcore_max_r == task_pcore_curr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:377:61  */
  assign n14314_o = n14313_o | task_lockstep_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:376:77  */
  assign n14315_o = n14314_o & n14312_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:376:15  */
  assign n14316_o = n14315_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:383:96  */
  assign delay_i_n14318 = delay_i_out_out; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:382:1  */
  delayv_16_1 delay_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(tid_rrrrrrrrrrr),
    .enable_in(n14319_o),
    .out_out(delay_i_out_out));
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14325_o = busy_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14326_o = ~n14325_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14327_o = delay_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14328_o = ~n14327_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14329_o = n14328_o & n14326_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14332_o = n14329_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14333_o = busy_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14334_o = ~n14333_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14335_o = delay_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14336_o = ~n14335_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14337_o = n14336_o & n14334_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14340_o = n14337_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14341_o = busy_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14342_o = ~n14341_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14343_o = delay_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14344_o = ~n14343_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14345_o = n14344_o & n14342_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14348_o = n14345_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14349_o = busy_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14350_o = ~n14349_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14351_o = delay_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14352_o = ~n14351_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14353_o = n14352_o & n14350_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14356_o = n14353_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14357_o = busy_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14358_o = ~n14357_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14359_o = delay_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14360_o = ~n14359_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14361_o = n14360_o & n14358_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14364_o = n14361_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14365_o = busy_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14366_o = ~n14365_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14367_o = delay_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14368_o = ~n14367_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14369_o = n14368_o & n14366_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14372_o = n14369_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14373_o = busy_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14374_o = ~n14373_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14375_o = delay_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14376_o = ~n14375_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14377_o = n14376_o & n14374_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14380_o = n14377_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14381_o = busy_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14382_o = ~n14381_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14383_o = delay_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14384_o = ~n14383_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14385_o = n14384_o & n14382_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14388_o = n14385_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14389_o = busy_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14390_o = ~n14389_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14391_o = delay_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14392_o = ~n14391_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14393_o = n14392_o & n14390_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14396_o = n14393_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14397_o = busy_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14398_o = ~n14397_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14399_o = delay_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14400_o = ~n14399_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14401_o = n14400_o & n14398_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14404_o = n14401_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14405_o = busy_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14406_o = ~n14405_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14407_o = delay_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14408_o = ~n14407_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14409_o = n14408_o & n14406_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14412_o = n14409_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14413_o = busy_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14414_o = ~n14413_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14415_o = delay_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14416_o = ~n14415_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14417_o = n14416_o & n14414_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14420_o = n14417_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14421_o = busy_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14422_o = ~n14421_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14423_o = delay_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14424_o = ~n14423_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14425_o = n14424_o & n14422_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14428_o = n14425_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14429_o = busy_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14430_o = ~n14429_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14431_o = delay_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14432_o = ~n14431_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14433_o = n14432_o & n14430_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14436_o = n14433_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14437_o = busy_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14438_o = ~n14437_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14439_o = delay_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14440_o = ~n14439_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14441_o = n14440_o & n14438_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14444_o = n14441_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:18  */
  assign n14445_o = busy_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:21  */
  assign n14446_o = ~n14445_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:37  */
  assign n14447_o = delay_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:394:40  */
  assign n14448_o = ~n14447_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:26  */
  assign n14449_o = n14448_o & n14446_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:394:9  */
  assign n14452_o = n14449_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14454_o = n14453_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14455_o = busy1[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14456_o = vm_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14457_o = ~n14456_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14458_o = n14455_o & n14457_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14459_o = n14454_o | n14458_o;
  assign n14461_o = n14460_o[1];
  assign n14462_o = {n14461_o, n14459_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14463_o = n14462_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14464_o = busy1[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14465_o = vm_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14466_o = n14464_o & n14465_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14467_o = n14463_o | n14466_o;
  assign n14468_o = {n14467_o, n14459_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14469_o = n14468_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14470_o = busy1[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14471_o = vm_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14472_o = ~n14471_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14473_o = n14470_o & n14472_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14474_o = n14469_o | n14473_o;
  assign n14475_o = {n14467_o, n14474_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14476_o = n14475_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14477_o = busy1[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14478_o = vm_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14479_o = n14477_o & n14478_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14480_o = n14476_o | n14479_o;
  assign n14481_o = {n14480_o, n14474_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14482_o = n14481_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14483_o = busy1[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14484_o = vm_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14485_o = ~n14484_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14486_o = n14483_o & n14485_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14487_o = n14482_o | n14486_o;
  assign n14488_o = {n14480_o, n14487_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14489_o = n14488_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14490_o = busy1[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14491_o = vm_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14492_o = n14490_o & n14491_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14493_o = n14489_o | n14492_o;
  assign n14494_o = {n14493_o, n14487_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14495_o = n14494_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14496_o = busy1[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14497_o = vm_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14498_o = ~n14497_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14499_o = n14496_o & n14498_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14500_o = n14495_o | n14499_o;
  assign n14501_o = {n14493_o, n14500_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14502_o = n14501_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14503_o = busy1[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14504_o = vm_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14505_o = n14503_o & n14504_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14506_o = n14502_o | n14505_o;
  assign n14507_o = {n14506_o, n14500_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14508_o = n14507_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14509_o = busy1[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14510_o = vm_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14511_o = ~n14510_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14512_o = n14509_o & n14511_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14513_o = n14508_o | n14512_o;
  assign n14514_o = {n14506_o, n14513_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14515_o = n14514_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14516_o = busy1[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14517_o = vm_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14518_o = n14516_o & n14517_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14519_o = n14515_o | n14518_o;
  assign n14520_o = {n14519_o, n14513_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14521_o = n14520_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14522_o = busy1[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14523_o = vm_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14524_o = ~n14523_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14525_o = n14522_o & n14524_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14526_o = n14521_o | n14525_o;
  assign n14527_o = {n14519_o, n14526_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14528_o = n14527_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14529_o = busy1[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14530_o = vm_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14531_o = n14529_o & n14530_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14532_o = n14528_o | n14531_o;
  assign n14533_o = {n14532_o, n14526_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14534_o = n14533_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14535_o = busy1[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14536_o = vm_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14537_o = ~n14536_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14538_o = n14535_o & n14537_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14539_o = n14534_o | n14538_o;
  assign n14540_o = {n14532_o, n14539_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14541_o = n14540_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14542_o = busy1[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14543_o = vm_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14544_o = n14542_o & n14543_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14545_o = n14541_o | n14544_o;
  assign n14546_o = {n14545_o, n14539_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14547_o = n14546_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14548_o = busy1[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14549_o = vm_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14550_o = ~n14549_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14551_o = n14548_o & n14550_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14552_o = n14547_o | n14551_o;
  assign n14553_o = {n14545_o, n14552_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14554_o = n14553_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14555_o = busy1[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14556_o = vm_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14557_o = n14555_o & n14556_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14558_o = n14554_o | n14557_o;
  assign n14559_o = {n14558_o, n14552_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14560_o = n14559_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14561_o = busy1[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14562_o = vm_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14563_o = ~n14562_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14564_o = n14561_o & n14563_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14565_o = n14560_o | n14564_o;
  assign n14566_o = {n14558_o, n14565_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14567_o = n14566_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14568_o = busy1[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14569_o = vm_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14570_o = n14568_o & n14569_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14571_o = n14567_o | n14570_o;
  assign n14572_o = {n14571_o, n14565_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14573_o = n14572_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14574_o = busy1[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14575_o = vm_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14576_o = ~n14575_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14577_o = n14574_o & n14576_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14578_o = n14573_o | n14577_o;
  assign n14579_o = {n14571_o, n14578_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14580_o = n14579_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14581_o = busy1[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14582_o = vm_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14583_o = n14581_o & n14582_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14584_o = n14580_o | n14583_o;
  assign n14585_o = {n14584_o, n14578_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14586_o = n14585_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14587_o = busy1[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14588_o = vm_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14589_o = ~n14588_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14590_o = n14587_o & n14589_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14591_o = n14586_o | n14590_o;
  assign n14592_o = {n14584_o, n14591_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14593_o = n14592_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14594_o = busy1[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14595_o = vm_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14596_o = n14594_o & n14595_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14597_o = n14593_o | n14596_o;
  assign n14598_o = {n14597_o, n14591_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14599_o = n14598_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14600_o = busy1[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14601_o = vm_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14602_o = ~n14601_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14603_o = n14600_o & n14602_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14604_o = n14599_o | n14603_o;
  assign n14605_o = {n14597_o, n14604_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14606_o = n14605_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14607_o = busy1[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14608_o = vm_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14609_o = n14607_o & n14608_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14610_o = n14606_o | n14609_o;
  assign n14611_o = {n14610_o, n14604_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14612_o = n14611_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14613_o = busy1[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14614_o = vm_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14615_o = ~n14614_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14616_o = n14613_o & n14615_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14617_o = n14612_o | n14616_o;
  assign n14618_o = {n14610_o, n14617_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14619_o = n14618_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14620_o = busy1[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14621_o = vm_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14622_o = n14620_o & n14621_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14623_o = n14619_o | n14622_o;
  assign n14624_o = {n14623_o, n14617_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14625_o = n14624_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14626_o = busy1[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14627_o = vm_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14628_o = ~n14627_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14629_o = n14626_o & n14628_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14630_o = n14625_o | n14629_o;
  assign n14631_o = {n14623_o, n14630_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14632_o = n14631_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14633_o = busy1[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14634_o = vm_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14635_o = n14633_o & n14634_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14636_o = n14632_o | n14635_o;
  assign n14637_o = {n14636_o, n14630_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14638_o = n14637_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14639_o = busy1[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14640_o = vm_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14641_o = ~n14640_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14642_o = n14639_o & n14641_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14643_o = n14638_o | n14642_o;
  assign n14644_o = {n14636_o, n14643_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14645_o = n14644_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14646_o = busy1[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14647_o = vm_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14648_o = n14646_o & n14647_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14649_o = n14645_o | n14648_o;
  assign n14650_o = {n14649_o, n14643_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:402:28  */
  assign n14651_o = n14650_o[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:41  */
  assign n14652_o = busy1[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:58  */
  assign n14653_o = vm_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:402:50  */
  assign n14654_o = ~n14653_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:45  */
  assign n14655_o = n14652_o & n14654_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:402:32  */
  assign n14656_o = n14651_o | n14655_o;
  assign n14657_o = {n14649_o, n14656_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:403:28  */
  assign n14658_o = n14657_o[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:41  */
  assign n14659_o = busy1[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:54  */
  assign n14660_o = vm_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:403:45  */
  assign n14661_o = n14659_o & n14660_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:403:32  */
  assign n14662_o = n14658_o | n14661_o;
  assign n14663_o = {n14662_o, n14656_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:414:16  */
  assign n14668_o = ~reset_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:450:51  */
  assign n14670_o = mu_instruction[79:75];
  /* ../../HW/src/pcore/instr_fetch.vhd:450:105  */
  assign n14672_o = n14670_o != 5'b00000;
  /* ../../HW/src/pcore/instr_fetch.vhd:450:33  */
  assign n14673_o = n14672_o & tid_valid_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:450:13  */
  assign n14676_o = n14673_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:455:54  */
  assign n14677_o = imu_instruction[31:27];
  /* ../../HW/src/pcore/instr_fetch.vhd:455:110  */
  assign n14679_o = n14677_o != 5'b00000;
  /* ../../HW/src/pcore/instr_fetch.vhd:455:35  */
  assign n14680_o = n14679_o & tid_valid_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:455:13  */
  assign n14683_o = n14680_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:280:11  */
  assign n14790_o = next_tid[7:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:280:24  */
  assign n14792_o = n14790_o == 8'b00000000;
  /* ../../HW/src/pcore/instr_fetch.vhd:281:14  */
  assign n14793_o = next_tid[11:8];
  /* ../../HW/src/pcore/instr_fetch.vhd:281:27  */
  assign n14795_o = n14793_o == 4'b0000;
  /* ../../HW/src/pcore/instr_fetch.vhd:282:17  */
  assign n14796_o = next_tid[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:284:20  */
  assign n14797_o = next_tid[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:286:20  */
  assign n14798_o = next_tid[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:286:11  */
  assign n14801_o = n14798_o ? 4'b1110 : 4'b1111;
  /* ../../HW/src/pcore/instr_fetch.vhd:284:11  */
  assign n14803_o = n14797_o ? 4'b1101 : n14801_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:282:11  */
  assign n14805_o = n14796_o ? 4'b1100 : n14803_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:292:17  */
  assign n14806_o = next_tid[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:294:20  */
  assign n14807_o = next_tid[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:296:20  */
  assign n14808_o = next_tid[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:296:11  */
  assign n14811_o = n14808_o ? 4'b1010 : 4'b1011;
  /* ../../HW/src/pcore/instr_fetch.vhd:294:11  */
  assign n14813_o = n14807_o ? 4'b1001 : n14811_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:292:11  */
  assign n14815_o = n14806_o ? 4'b1000 : n14813_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:281:8  */
  assign n14816_o = n14795_o ? n14805_o : n14815_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:303:14  */
  assign n14817_o = next_tid[3:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:303:26  */
  assign n14819_o = n14817_o == 4'b0000;
  /* ../../HW/src/pcore/instr_fetch.vhd:304:17  */
  assign n14820_o = next_tid[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:306:20  */
  assign n14821_o = next_tid[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:308:20  */
  assign n14822_o = next_tid[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:308:11  */
  assign n14825_o = n14822_o ? 4'b0110 : 4'b0111;
  /* ../../HW/src/pcore/instr_fetch.vhd:306:11  */
  assign n14827_o = n14821_o ? 4'b0101 : n14825_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:304:11  */
  assign n14829_o = n14820_o ? 4'b0100 : n14827_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:314:17  */
  assign n14830_o = next_tid[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:316:20  */
  assign n14831_o = next_tid[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:318:20  */
  assign n14832_o = next_tid[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:318:11  */
  assign n14835_o = n14832_o ? 4'b0010 : 4'b0011;
  /* ../../HW/src/pcore/instr_fetch.vhd:316:11  */
  assign n14837_o = n14831_o ? 4'b0001 : n14835_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:314:11  */
  assign n14839_o = n14830_o ? 4'b0000 : n14837_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:303:8  */
  assign n14840_o = n14819_o ? n14829_o : n14839_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:280:5  */
  assign n14841_o = n14792_o ? n14816_o : n14840_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:512:34  */
  assign arbiter_1_i_n14843 = arbiter_1_i_gnt_out; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:513:40  */
  assign arbiter_1_i_n14844 = arbiter_1_i_gnt_valid_out; // (signal)
  /* ../../HW/src/pcore/instr_fetch.vhd:504:1  */
  arbiter_16_5ba93c9db0cff93f52b521d7420e43f6eda2784f arbiter_1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .req_in(avail),
    .gnt_out(arbiter_1_i_gnt_out),
    .gnt_valid_out(arbiter_1_i_gnt_valid_out));
  /* ../../HW/src/pcore/instr_fetch.vhd:520:20  */
  assign n14849_o = tid_rrrrrrr | tid_rrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:520:34  */
  assign n14850_o = n14849_o | tid_rrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:520:47  */
  assign n14851_o = n14850_o | tid_rrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:520:59  */
  assign n14852_o = n14851_o | tid_rrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:520:70  */
  assign n14853_o = n14852_o | tid_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:520:80  */
  assign n14854_o = n14853_o | tid_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:254:4  */
  assign n14862_o = task_tid_mask_in == 4'b0000;
  /* ../../HW/src/pcore/instr_fetch.vhd:255:4  */
  assign n14864_o = task_tid_mask_in == 4'b0001;
  /* ../../HW/src/pcore/instr_fetch.vhd:256:4  */
  assign n14866_o = task_tid_mask_in == 4'b0010;
  /* ../../HW/src/pcore/instr_fetch.vhd:257:4  */
  assign n14868_o = task_tid_mask_in == 4'b0011;
  /* ../../HW/src/pcore/instr_fetch.vhd:258:4  */
  assign n14870_o = task_tid_mask_in == 4'b0100;
  /* ../../HW/src/pcore/instr_fetch.vhd:259:4  */
  assign n14872_o = task_tid_mask_in == 4'b0101;
  /* ../../HW/src/pcore/instr_fetch.vhd:260:4  */
  assign n14874_o = task_tid_mask_in == 4'b0110;
  /* ../../HW/src/pcore/instr_fetch.vhd:261:4  */
  assign n14876_o = task_tid_mask_in == 4'b0111;
  /* ../../HW/src/pcore/instr_fetch.vhd:262:4  */
  assign n14878_o = task_tid_mask_in == 4'b1000;
  /* ../../HW/src/pcore/instr_fetch.vhd:263:4  */
  assign n14880_o = task_tid_mask_in == 4'b1001;
  /* ../../HW/src/pcore/instr_fetch.vhd:264:4  */
  assign n14882_o = task_tid_mask_in == 4'b1010;
  /* ../../HW/src/pcore/instr_fetch.vhd:265:4  */
  assign n14884_o = task_tid_mask_in == 4'b1011;
  /* ../../HW/src/pcore/instr_fetch.vhd:266:4  */
  assign n14886_o = task_tid_mask_in == 4'b1100;
  /* ../../HW/src/pcore/instr_fetch.vhd:267:4  */
  assign n14888_o = task_tid_mask_in == 4'b1101;
  /* ../../HW/src/pcore/instr_fetch.vhd:268:4  */
  assign n14890_o = task_tid_mask_in == 4'b1110;
  assign n14891_o = {n14890_o, n14888_o, n14886_o, n14884_o, n14882_o, n14880_o, n14878_o, n14876_o, n14874_o, n14872_o, n14870_o, n14868_o, n14866_o, n14864_o, n14862_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:253:1  */
  always @*
    case (n14891_o)
      15'b100000000000000: n14908_o = 16'b0111111111111111;
      15'b010000000000000: n14908_o = 16'b0011111111111111;
      15'b001000000000000: n14908_o = 16'b0001111111111111;
      15'b000100000000000: n14908_o = 16'b0000111111111111;
      15'b000010000000000: n14908_o = 16'b0000011111111111;
      15'b000001000000000: n14908_o = 16'b0000001111111111;
      15'b000000100000000: n14908_o = 16'b0000000111111111;
      15'b000000010000000: n14908_o = 16'b0000000011111111;
      15'b000000001000000: n14908_o = 16'b0000000001111111;
      15'b000000000100000: n14908_o = 16'b0000000000111111;
      15'b000000000010000: n14908_o = 16'b0000000000011111;
      15'b000000000001000: n14908_o = 16'b0000000000001111;
      15'b000000000000100: n14908_o = 16'b0000000000000111;
      15'b000000000000010: n14908_o = 16'b0000000000000011;
      15'b000000000000001: n14908_o = 16'b0000000000000001;
      default: n14908_o = 16'b1111111111111111;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:536:16  */
  assign n14918_o = ~reset_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n14923_o = task_in ? 5'b00000 : task_pcore_curr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:23  */
  assign n14931_o = task_mask_r == 16'b0000000000000000;
  /* ../../HW/src/pcore/instr_fetch.vhd:584:29  */
  assign n14932_o = task_pcore_max_r != task_pcore_curr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:67  */
  assign n14933_o = n14932_o & n14931_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:585:26  */
  assign n14934_o = ~task_lockstep_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:584:51  */
  assign n14935_o = n14934_o & n14933_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:586:17  */
  assign n14937_o = busy_r == 16'b0000000000000000;
  /* ../../HW/src/pcore/instr_fetch.vhd:585:31  */
  assign n14938_o = n14937_o & n14935_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:587:59  */
  assign n14940_o = task_pcore_curr_r + 5'b00001;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n14941_o = n14938_o ? n14940_o : n14923_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n14943_o = busy_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n14944_o = ~n14943_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n14945_o = task_mask_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n14946_o = n14945_o & n14944_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n14947_o = tid_rrrrrrrrrrr[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n14948_o = ~n14947_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n14949_o = n14948_o & n14946_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n14951_o = tid[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n14952_o = tid_delay[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n14953_o = delay_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n14955_o = n14952_o ? 1'b0 : n14953_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n14957_o = n14951_o ? 1'b1 : n14955_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n14958_o = vm_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n14959_o = data_model_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n14960_o = tid_rrrrrrrrrrr[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n14961_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n14962_o = pc_r[175:165];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n14963_o = busy_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n14964_o = tid[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n14965_o = tid_delay[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n14966_o = delay_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n14968_o = n14965_o ? 1'b0 : n14966_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n14970_o = n14964_o ? 1'b1 : n14968_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n14971_o = n14960_o ? next_addr : n14962_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n14972_o = n14960_o ? n14961_o : n14963_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n14974_o = n14960_o ? 1'b1 : n14970_o;
  assign n14975_o = task_tid_mask_r[0];
  assign n14976_o = task_tid_mask[0];
  assign n14977_o = task_mask_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n14978_o = task_in ? n14976_o : n14977_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n14979_o = n14938_o ? n14975_o : n14978_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14980_o = n14949_o ? 1'b0 : n14979_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14986_o = n14949_o ? task_start_addr_r : n14971_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14988_o = n14949_o ? 1'b1 : n14972_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14989_o = n14949_o ? n14957_o : n14974_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14990_o = n14949_o ? task_vm_r : n14958_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14991_o = n14949_o ? task2_data_model_r : n14959_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n14994_o = n14949_o ? 1'b1 : 1'b0;
  assign n14995_o = iregister_auto_r[27:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n14996_o = n14994_o ? task_iregister_auto_r : n14995_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n14997_o = ~n14989_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n14998_o = n14997_o & n14988_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n14999_o = next_tid[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15000_o = ~n14999_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15001_o = n15000_o & n14998_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15004_o = n15001_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15005_o = busy_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15006_o = ~n15005_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15007_o = task_mask_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15008_o = n15007_o & n15006_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15009_o = tid_rrrrrrrrrrr[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15010_o = ~n15009_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15011_o = n15010_o & n15008_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15013_o = tid[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15014_o = tid_delay[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15015_o = delay_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15017_o = n15014_o ? 1'b0 : n15015_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15019_o = n15013_o ? 1'b1 : n15017_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15020_o = vm_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15021_o = data_model_r[3:2];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15022_o = tid_rrrrrrrrrrr[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15023_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15024_o = pc_r[164:154];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15025_o = busy_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15026_o = tid[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15027_o = tid_delay[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15028_o = delay_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15030_o = n15027_o ? 1'b0 : n15028_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15032_o = n15026_o ? 1'b1 : n15030_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15033_o = n15022_o ? next_addr : n15024_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15034_o = n15022_o ? n15023_o : n15025_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15036_o = n15022_o ? 1'b1 : n15032_o;
  assign n15037_o = task_tid_mask_r[1];
  assign n15038_o = task_tid_mask[1];
  assign n15039_o = task_mask_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15040_o = task_in ? n15038_o : n15039_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15041_o = n14938_o ? n15037_o : n15040_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15042_o = n15011_o ? 1'b0 : n15041_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15048_o = n15011_o ? task_start_addr_r : n15033_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15050_o = n15011_o ? 1'b1 : n15034_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15051_o = n15011_o ? n15019_o : n15036_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15052_o = n15011_o ? task_vm_r : n15020_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15053_o = n15011_o ? task2_data_model_r : n15021_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15056_o = n15011_o ? 1'b1 : 1'b0;
  assign n15057_o = iregister_auto_r[55:28];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15058_o = n15056_o ? task_iregister_auto_r : n15057_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15059_o = ~n15051_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15060_o = n15059_o & n15050_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15061_o = next_tid[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15062_o = ~n15061_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15063_o = n15062_o & n15060_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15066_o = n15063_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15067_o = busy_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15068_o = ~n15067_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15069_o = task_mask_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15070_o = n15069_o & n15068_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15071_o = tid_rrrrrrrrrrr[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15072_o = ~n15071_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15073_o = n15072_o & n15070_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15075_o = tid[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15076_o = tid_delay[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15077_o = delay_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15079_o = n15076_o ? 1'b0 : n15077_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15081_o = n15075_o ? 1'b1 : n15079_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15082_o = vm_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15083_o = data_model_r[5:4];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15084_o = tid_rrrrrrrrrrr[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15085_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15086_o = pc_r[153:143];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15087_o = busy_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15088_o = tid[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15089_o = tid_delay[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15090_o = delay_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15092_o = n15089_o ? 1'b0 : n15090_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15094_o = n15088_o ? 1'b1 : n15092_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15095_o = n15084_o ? next_addr : n15086_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15096_o = n15084_o ? n15085_o : n15087_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15098_o = n15084_o ? 1'b1 : n15094_o;
  assign n15099_o = task_tid_mask_r[2];
  assign n15100_o = task_tid_mask[2];
  assign n15101_o = task_mask_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15102_o = task_in ? n15100_o : n15101_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15103_o = n14938_o ? n15099_o : n15102_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15104_o = n15073_o ? 1'b0 : n15103_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15110_o = n15073_o ? task_start_addr_r : n15095_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15112_o = n15073_o ? 1'b1 : n15096_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15113_o = n15073_o ? n15081_o : n15098_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15114_o = n15073_o ? task_vm_r : n15082_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15115_o = n15073_o ? task2_data_model_r : n15083_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15118_o = n15073_o ? 1'b1 : 1'b0;
  assign n15119_o = iregister_auto_r[83:56];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15120_o = n15118_o ? task_iregister_auto_r : n15119_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15121_o = ~n15113_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15122_o = n15121_o & n15112_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15123_o = next_tid[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15124_o = ~n15123_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15125_o = n15124_o & n15122_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15128_o = n15125_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15129_o = busy_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15130_o = ~n15129_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15131_o = task_mask_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15132_o = n15131_o & n15130_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15133_o = tid_rrrrrrrrrrr[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15134_o = ~n15133_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15135_o = n15134_o & n15132_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15137_o = tid[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15138_o = tid_delay[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15139_o = delay_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15141_o = n15138_o ? 1'b0 : n15139_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15143_o = n15137_o ? 1'b1 : n15141_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15144_o = vm_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15145_o = data_model_r[7:6];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15146_o = tid_rrrrrrrrrrr[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15147_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15148_o = pc_r[142:132];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15149_o = busy_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15150_o = tid[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15151_o = tid_delay[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15152_o = delay_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15154_o = n15151_o ? 1'b0 : n15152_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15156_o = n15150_o ? 1'b1 : n15154_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15157_o = n15146_o ? next_addr : n15148_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15158_o = n15146_o ? n15147_o : n15149_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15160_o = n15146_o ? 1'b1 : n15156_o;
  assign n15161_o = task_tid_mask_r[3];
  assign n15162_o = task_tid_mask[3];
  assign n15163_o = task_mask_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15164_o = task_in ? n15162_o : n15163_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15165_o = n14938_o ? n15161_o : n15164_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15166_o = n15135_o ? 1'b0 : n15165_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15172_o = n15135_o ? task_start_addr_r : n15157_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15174_o = n15135_o ? 1'b1 : n15158_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15175_o = n15135_o ? n15143_o : n15160_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15176_o = n15135_o ? task_vm_r : n15144_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15177_o = n15135_o ? task2_data_model_r : n15145_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15180_o = n15135_o ? 1'b1 : 1'b0;
  assign n15181_o = iregister_auto_r[111:84];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15182_o = n15180_o ? task_iregister_auto_r : n15181_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15183_o = ~n15175_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15184_o = n15183_o & n15174_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15185_o = next_tid[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15186_o = ~n15185_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15187_o = n15186_o & n15184_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15190_o = n15187_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15191_o = busy_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15192_o = ~n15191_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15193_o = task_mask_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15194_o = n15193_o & n15192_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15195_o = tid_rrrrrrrrrrr[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15196_o = ~n15195_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15197_o = n15196_o & n15194_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15199_o = tid[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15200_o = tid_delay[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15201_o = delay_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15203_o = n15200_o ? 1'b0 : n15201_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15205_o = n15199_o ? 1'b1 : n15203_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15206_o = vm_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15207_o = data_model_r[9:8];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15208_o = tid_rrrrrrrrrrr[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15209_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15210_o = pc_r[131:121];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15211_o = busy_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15212_o = tid[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15213_o = tid_delay[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15214_o = delay_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15216_o = n15213_o ? 1'b0 : n15214_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15218_o = n15212_o ? 1'b1 : n15216_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15219_o = n15208_o ? next_addr : n15210_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15220_o = n15208_o ? n15209_o : n15211_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15222_o = n15208_o ? 1'b1 : n15218_o;
  assign n15223_o = task_tid_mask_r[4];
  assign n15224_o = task_tid_mask[4];
  assign n15225_o = task_mask_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15226_o = task_in ? n15224_o : n15225_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15227_o = n14938_o ? n15223_o : n15226_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15228_o = n15197_o ? 1'b0 : n15227_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15234_o = n15197_o ? task_start_addr_r : n15219_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15236_o = n15197_o ? 1'b1 : n15220_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15237_o = n15197_o ? n15205_o : n15222_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15238_o = n15197_o ? task_vm_r : n15206_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15239_o = n15197_o ? task2_data_model_r : n15207_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15242_o = n15197_o ? 1'b1 : 1'b0;
  assign n15243_o = iregister_auto_r[139:112];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15244_o = n15242_o ? task_iregister_auto_r : n15243_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15245_o = ~n15237_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15246_o = n15245_o & n15236_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15247_o = next_tid[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15248_o = ~n15247_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15249_o = n15248_o & n15246_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15252_o = n15249_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15253_o = busy_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15254_o = ~n15253_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15255_o = task_mask_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15256_o = n15255_o & n15254_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15257_o = tid_rrrrrrrrrrr[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15258_o = ~n15257_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15259_o = n15258_o & n15256_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15261_o = tid[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15262_o = tid_delay[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15263_o = delay_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15265_o = n15262_o ? 1'b0 : n15263_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15267_o = n15261_o ? 1'b1 : n15265_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15268_o = vm_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15269_o = data_model_r[11:10];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15270_o = tid_rrrrrrrrrrr[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15271_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15272_o = pc_r[120:110];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15273_o = busy_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15274_o = tid[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15275_o = tid_delay[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15276_o = delay_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15278_o = n15275_o ? 1'b0 : n15276_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15280_o = n15274_o ? 1'b1 : n15278_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15281_o = n15270_o ? next_addr : n15272_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15282_o = n15270_o ? n15271_o : n15273_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15284_o = n15270_o ? 1'b1 : n15280_o;
  assign n15285_o = task_tid_mask_r[5];
  assign n15286_o = task_tid_mask[5];
  assign n15287_o = task_mask_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15288_o = task_in ? n15286_o : n15287_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15289_o = n14938_o ? n15285_o : n15288_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15290_o = n15259_o ? 1'b0 : n15289_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15296_o = n15259_o ? task_start_addr_r : n15281_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15298_o = n15259_o ? 1'b1 : n15282_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15299_o = n15259_o ? n15267_o : n15284_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15300_o = n15259_o ? task_vm_r : n15268_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15301_o = n15259_o ? task2_data_model_r : n15269_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15304_o = n15259_o ? 1'b1 : 1'b0;
  assign n15305_o = iregister_auto_r[167:140];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15306_o = n15304_o ? task_iregister_auto_r : n15305_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15307_o = ~n15299_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15308_o = n15307_o & n15298_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15309_o = next_tid[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15310_o = ~n15309_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15311_o = n15310_o & n15308_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15314_o = n15311_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15315_o = busy_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15316_o = ~n15315_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15317_o = task_mask_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15318_o = n15317_o & n15316_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15319_o = tid_rrrrrrrrrrr[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15320_o = ~n15319_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15321_o = n15320_o & n15318_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15323_o = tid[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15324_o = tid_delay[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15325_o = delay_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15327_o = n15324_o ? 1'b0 : n15325_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15329_o = n15323_o ? 1'b1 : n15327_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15330_o = vm_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15331_o = data_model_r[13:12];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15332_o = tid_rrrrrrrrrrr[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15333_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15334_o = pc_r[109:99];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15335_o = busy_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15336_o = tid[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15337_o = tid_delay[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15338_o = delay_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15340_o = n15337_o ? 1'b0 : n15338_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15342_o = n15336_o ? 1'b1 : n15340_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15343_o = n15332_o ? next_addr : n15334_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15344_o = n15332_o ? n15333_o : n15335_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15346_o = n15332_o ? 1'b1 : n15342_o;
  assign n15347_o = task_tid_mask_r[6];
  assign n15348_o = task_tid_mask[6];
  assign n15349_o = task_mask_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15350_o = task_in ? n15348_o : n15349_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15351_o = n14938_o ? n15347_o : n15350_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15352_o = n15321_o ? 1'b0 : n15351_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15358_o = n15321_o ? task_start_addr_r : n15343_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15360_o = n15321_o ? 1'b1 : n15344_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15361_o = n15321_o ? n15329_o : n15346_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15362_o = n15321_o ? task_vm_r : n15330_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15363_o = n15321_o ? task2_data_model_r : n15331_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15366_o = n15321_o ? 1'b1 : 1'b0;
  assign n15367_o = iregister_auto_r[195:168];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15368_o = n15366_o ? task_iregister_auto_r : n15367_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15369_o = ~n15361_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15370_o = n15369_o & n15360_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15371_o = next_tid[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15372_o = ~n15371_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15373_o = n15372_o & n15370_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15376_o = n15373_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15377_o = busy_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15378_o = ~n15377_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15379_o = task_mask_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15380_o = n15379_o & n15378_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15381_o = tid_rrrrrrrrrrr[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15382_o = ~n15381_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15383_o = n15382_o & n15380_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15385_o = tid[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15386_o = tid_delay[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15387_o = delay_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15389_o = n15386_o ? 1'b0 : n15387_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15391_o = n15385_o ? 1'b1 : n15389_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15392_o = vm_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15393_o = data_model_r[15:14];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15394_o = tid_rrrrrrrrrrr[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15395_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15396_o = pc_r[98:88];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15397_o = busy_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15398_o = tid[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15399_o = tid_delay[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15400_o = delay_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15402_o = n15399_o ? 1'b0 : n15400_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15404_o = n15398_o ? 1'b1 : n15402_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15405_o = n15394_o ? next_addr : n15396_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15406_o = n15394_o ? n15395_o : n15397_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15408_o = n15394_o ? 1'b1 : n15404_o;
  assign n15409_o = task_tid_mask_r[7];
  assign n15410_o = task_tid_mask[7];
  assign n15411_o = task_mask_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15412_o = task_in ? n15410_o : n15411_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15413_o = n14938_o ? n15409_o : n15412_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15414_o = n15383_o ? 1'b0 : n15413_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15420_o = n15383_o ? task_start_addr_r : n15405_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15422_o = n15383_o ? 1'b1 : n15406_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15423_o = n15383_o ? n15391_o : n15408_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15424_o = n15383_o ? task_vm_r : n15392_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15425_o = n15383_o ? task2_data_model_r : n15393_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15428_o = n15383_o ? 1'b1 : 1'b0;
  assign n15429_o = iregister_auto_r[223:196];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15430_o = n15428_o ? task_iregister_auto_r : n15429_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15431_o = ~n15423_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15432_o = n15431_o & n15422_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15433_o = next_tid[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15434_o = ~n15433_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15435_o = n15434_o & n15432_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15438_o = n15435_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15439_o = busy_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15440_o = ~n15439_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15441_o = task_mask_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15442_o = n15441_o & n15440_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15443_o = tid_rrrrrrrrrrr[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15444_o = ~n15443_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15445_o = n15444_o & n15442_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15447_o = tid[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15448_o = tid_delay[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15449_o = delay_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15451_o = n15448_o ? 1'b0 : n15449_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15453_o = n15447_o ? 1'b1 : n15451_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15454_o = vm_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15455_o = data_model_r[17:16];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15456_o = tid_rrrrrrrrrrr[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15457_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15458_o = pc_r[87:77];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15459_o = busy_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15460_o = tid[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15461_o = tid_delay[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15462_o = delay_r[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15464_o = n15461_o ? 1'b0 : n15462_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15466_o = n15460_o ? 1'b1 : n15464_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15467_o = n15456_o ? next_addr : n15458_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15468_o = n15456_o ? n15457_o : n15459_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15470_o = n15456_o ? 1'b1 : n15466_o;
  assign n15471_o = task_tid_mask_r[8];
  assign n15472_o = task_tid_mask[8];
  assign n15473_o = task_mask_r[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15474_o = task_in ? n15472_o : n15473_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15475_o = n14938_o ? n15471_o : n15474_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15476_o = n15445_o ? 1'b0 : n15475_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15482_o = n15445_o ? task_start_addr_r : n15467_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15484_o = n15445_o ? 1'b1 : n15468_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15485_o = n15445_o ? n15453_o : n15470_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15486_o = n15445_o ? task_vm_r : n15454_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15487_o = n15445_o ? task2_data_model_r : n15455_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15490_o = n15445_o ? 1'b1 : 1'b0;
  assign n15491_o = iregister_auto_r[251:224];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15492_o = n15490_o ? task_iregister_auto_r : n15491_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15493_o = ~n15485_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15494_o = n15493_o & n15484_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15495_o = next_tid[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15496_o = ~n15495_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15497_o = n15496_o & n15494_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15500_o = n15497_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15501_o = busy_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15502_o = ~n15501_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15503_o = task_mask_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15504_o = n15503_o & n15502_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15505_o = tid_rrrrrrrrrrr[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15506_o = ~n15505_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15507_o = n15506_o & n15504_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15509_o = tid[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15510_o = tid_delay[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15511_o = delay_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15513_o = n15510_o ? 1'b0 : n15511_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15515_o = n15509_o ? 1'b1 : n15513_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15516_o = vm_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15517_o = data_model_r[19:18];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15518_o = tid_rrrrrrrrrrr[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15519_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15520_o = pc_r[76:66];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15521_o = busy_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15522_o = tid[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15523_o = tid_delay[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15524_o = delay_r[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15526_o = n15523_o ? 1'b0 : n15524_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15528_o = n15522_o ? 1'b1 : n15526_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15529_o = n15518_o ? next_addr : n15520_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15530_o = n15518_o ? n15519_o : n15521_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15532_o = n15518_o ? 1'b1 : n15528_o;
  assign n15533_o = task_tid_mask_r[9];
  assign n15534_o = task_tid_mask[9];
  assign n15535_o = task_mask_r[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15536_o = task_in ? n15534_o : n15535_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15537_o = n14938_o ? n15533_o : n15536_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15538_o = n15507_o ? 1'b0 : n15537_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15544_o = n15507_o ? task_start_addr_r : n15529_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15546_o = n15507_o ? 1'b1 : n15530_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15547_o = n15507_o ? n15515_o : n15532_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15548_o = n15507_o ? task_vm_r : n15516_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15549_o = n15507_o ? task2_data_model_r : n15517_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15552_o = n15507_o ? 1'b1 : 1'b0;
  assign n15553_o = iregister_auto_r[279:252];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15554_o = n15552_o ? task_iregister_auto_r : n15553_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15555_o = ~n15547_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15556_o = n15555_o & n15546_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15557_o = next_tid[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15558_o = ~n15557_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15559_o = n15558_o & n15556_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15562_o = n15559_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15563_o = busy_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15564_o = ~n15563_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15565_o = task_mask_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15566_o = n15565_o & n15564_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15567_o = tid_rrrrrrrrrrr[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15568_o = ~n15567_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15569_o = n15568_o & n15566_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15571_o = tid[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15572_o = tid_delay[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15573_o = delay_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15575_o = n15572_o ? 1'b0 : n15573_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15577_o = n15571_o ? 1'b1 : n15575_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15578_o = vm_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15579_o = data_model_r[21:20];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15580_o = tid_rrrrrrrrrrr[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15581_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15582_o = pc_r[65:55];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15583_o = busy_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15584_o = tid[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15585_o = tid_delay[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15586_o = delay_r[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15588_o = n15585_o ? 1'b0 : n15586_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15590_o = n15584_o ? 1'b1 : n15588_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15591_o = n15580_o ? next_addr : n15582_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15592_o = n15580_o ? n15581_o : n15583_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15594_o = n15580_o ? 1'b1 : n15590_o;
  assign n15595_o = task_tid_mask_r[10];
  assign n15596_o = task_tid_mask[10];
  assign n15597_o = task_mask_r[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15598_o = task_in ? n15596_o : n15597_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15599_o = n14938_o ? n15595_o : n15598_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15600_o = n15569_o ? 1'b0 : n15599_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15606_o = n15569_o ? task_start_addr_r : n15591_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15608_o = n15569_o ? 1'b1 : n15592_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15609_o = n15569_o ? n15577_o : n15594_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15610_o = n15569_o ? task_vm_r : n15578_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15611_o = n15569_o ? task2_data_model_r : n15579_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15614_o = n15569_o ? 1'b1 : 1'b0;
  assign n15615_o = iregister_auto_r[307:280];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15616_o = n15614_o ? task_iregister_auto_r : n15615_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15617_o = ~n15609_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15618_o = n15617_o & n15608_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15619_o = next_tid[10];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15620_o = ~n15619_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15621_o = n15620_o & n15618_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15624_o = n15621_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15625_o = busy_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15626_o = ~n15625_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15627_o = task_mask_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15628_o = n15627_o & n15626_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15629_o = tid_rrrrrrrrrrr[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15630_o = ~n15629_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15631_o = n15630_o & n15628_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15633_o = tid[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15634_o = tid_delay[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15635_o = delay_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15637_o = n15634_o ? 1'b0 : n15635_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15639_o = n15633_o ? 1'b1 : n15637_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15640_o = vm_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15641_o = data_model_r[23:22];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15642_o = tid_rrrrrrrrrrr[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15643_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15644_o = pc_r[54:44];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15645_o = busy_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15646_o = tid[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15647_o = tid_delay[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15648_o = delay_r[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15650_o = n15647_o ? 1'b0 : n15648_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15652_o = n15646_o ? 1'b1 : n15650_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15653_o = n15642_o ? next_addr : n15644_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15654_o = n15642_o ? n15643_o : n15645_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15656_o = n15642_o ? 1'b1 : n15652_o;
  assign n15657_o = task_tid_mask_r[11];
  assign n15658_o = task_tid_mask[11];
  assign n15659_o = task_mask_r[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15660_o = task_in ? n15658_o : n15659_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15661_o = n14938_o ? n15657_o : n15660_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15662_o = n15631_o ? 1'b0 : n15661_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15668_o = n15631_o ? task_start_addr_r : n15653_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15670_o = n15631_o ? 1'b1 : n15654_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15671_o = n15631_o ? n15639_o : n15656_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15672_o = n15631_o ? task_vm_r : n15640_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15673_o = n15631_o ? task2_data_model_r : n15641_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15676_o = n15631_o ? 1'b1 : 1'b0;
  assign n15677_o = iregister_auto_r[335:308];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15678_o = n15676_o ? task_iregister_auto_r : n15677_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15679_o = ~n15671_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15680_o = n15679_o & n15670_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15681_o = next_tid[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15682_o = ~n15681_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15683_o = n15682_o & n15680_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15686_o = n15683_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15687_o = busy_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15688_o = ~n15687_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15689_o = task_mask_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15690_o = n15689_o & n15688_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15691_o = tid_rrrrrrrrrrr[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15692_o = ~n15691_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15693_o = n15692_o & n15690_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15695_o = tid[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15696_o = tid_delay[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15697_o = delay_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15699_o = n15696_o ? 1'b0 : n15697_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15701_o = n15695_o ? 1'b1 : n15699_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15702_o = vm_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15703_o = data_model_r[25:24];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15704_o = tid_rrrrrrrrrrr[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15705_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15706_o = pc_r[43:33];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15707_o = busy_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15708_o = tid[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15709_o = tid_delay[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15710_o = delay_r[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15712_o = n15709_o ? 1'b0 : n15710_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15714_o = n15708_o ? 1'b1 : n15712_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15715_o = n15704_o ? next_addr : n15706_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15716_o = n15704_o ? n15705_o : n15707_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15718_o = n15704_o ? 1'b1 : n15714_o;
  assign n15719_o = task_tid_mask_r[12];
  assign n15720_o = task_tid_mask[12];
  assign n15721_o = task_mask_r[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15722_o = task_in ? n15720_o : n15721_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15723_o = n14938_o ? n15719_o : n15722_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15724_o = n15693_o ? 1'b0 : n15723_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15730_o = n15693_o ? task_start_addr_r : n15715_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15732_o = n15693_o ? 1'b1 : n15716_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15733_o = n15693_o ? n15701_o : n15718_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15734_o = n15693_o ? task_vm_r : n15702_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15735_o = n15693_o ? task2_data_model_r : n15703_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15738_o = n15693_o ? 1'b1 : 1'b0;
  assign n15739_o = iregister_auto_r[363:336];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15740_o = n15738_o ? task_iregister_auto_r : n15739_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15741_o = ~n15733_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15742_o = n15741_o & n15732_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15743_o = next_tid[12];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15744_o = ~n15743_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15745_o = n15744_o & n15742_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15748_o = n15745_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15749_o = busy_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15750_o = ~n15749_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15751_o = task_mask_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15752_o = n15751_o & n15750_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15753_o = tid_rrrrrrrrrrr[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15754_o = ~n15753_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15755_o = n15754_o & n15752_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15757_o = tid[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15758_o = tid_delay[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15759_o = delay_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15761_o = n15758_o ? 1'b0 : n15759_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15763_o = n15757_o ? 1'b1 : n15761_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15764_o = vm_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15765_o = data_model_r[27:26];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15766_o = tid_rrrrrrrrrrr[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15767_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15768_o = pc_r[32:22];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15769_o = busy_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15770_o = tid[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15771_o = tid_delay[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15772_o = delay_r[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15774_o = n15771_o ? 1'b0 : n15772_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15776_o = n15770_o ? 1'b1 : n15774_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15777_o = n15766_o ? next_addr : n15768_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15778_o = n15766_o ? n15767_o : n15769_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15780_o = n15766_o ? 1'b1 : n15776_o;
  assign n15781_o = task_tid_mask_r[13];
  assign n15782_o = task_tid_mask[13];
  assign n15783_o = task_mask_r[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15784_o = task_in ? n15782_o : n15783_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15785_o = n14938_o ? n15781_o : n15784_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15786_o = n15755_o ? 1'b0 : n15785_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15792_o = n15755_o ? task_start_addr_r : n15777_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15794_o = n15755_o ? 1'b1 : n15778_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15795_o = n15755_o ? n15763_o : n15780_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15796_o = n15755_o ? task_vm_r : n15764_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15797_o = n15755_o ? task2_data_model_r : n15765_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15800_o = n15755_o ? 1'b1 : 1'b0;
  assign n15801_o = iregister_auto_r[391:364];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15802_o = n15800_o ? task_iregister_auto_r : n15801_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15803_o = ~n15795_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15804_o = n15803_o & n15794_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15805_o = next_tid[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15806_o = ~n15805_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15807_o = n15806_o & n15804_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15810_o = n15807_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15811_o = busy_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15812_o = ~n15811_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15813_o = task_mask_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15814_o = n15813_o & n15812_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15815_o = tid_rrrrrrrrrrr[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15816_o = ~n15815_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15817_o = n15816_o & n15814_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15819_o = tid[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15820_o = tid_delay[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15821_o = delay_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15823_o = n15820_o ? 1'b0 : n15821_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15825_o = n15819_o ? 1'b1 : n15823_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15826_o = vm_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15827_o = data_model_r[29:28];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15828_o = tid_rrrrrrrrrrr[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15829_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15830_o = pc_r[21:11];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15831_o = busy_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15832_o = tid[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15833_o = tid_delay[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15834_o = delay_r[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15836_o = n15833_o ? 1'b0 : n15834_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15838_o = n15832_o ? 1'b1 : n15836_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15839_o = n15828_o ? next_addr : n15830_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15840_o = n15828_o ? n15829_o : n15831_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15842_o = n15828_o ? 1'b1 : n15838_o;
  assign n15843_o = task_tid_mask_r[14];
  assign n15844_o = task_tid_mask[14];
  assign n15845_o = task_mask_r[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15846_o = task_in ? n15844_o : n15845_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15847_o = n14938_o ? n15843_o : n15846_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15848_o = n15817_o ? 1'b0 : n15847_o;
  assign n15849_o = task_tid_mask_r[15];
  assign n15850_o = task_tid_mask[15];
  assign n15851_o = task_mask_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n15852_o = task_in ? n15850_o : n15851_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n15853_o = n14938_o ? n15849_o : n15852_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15854_o = n15817_o ? task_start_addr_r : n15839_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15856_o = n15817_o ? 1'b1 : n15840_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15857_o = n15817_o ? n15825_o : n15842_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15858_o = n15817_o ? task_vm_r : n15826_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15859_o = n15817_o ? task2_data_model_r : n15827_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15862_o = n15817_o ? 1'b1 : 1'b0;
  assign n15863_o = iregister_auto_r[419:392];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15864_o = n15862_o ? task_iregister_auto_r : n15863_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15865_o = ~n15857_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15866_o = n15865_o & n15856_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15867_o = next_tid[14];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15868_o = ~n15867_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15869_o = n15868_o & n15866_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15872_o = n15869_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:21  */
  assign n15873_o = busy_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:24  */
  assign n15874_o = ~n15873_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:44  */
  assign n15875_o = task_mask_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:29  */
  assign n15876_o = n15875_o & n15874_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:71  */
  assign n15877_o = tid_rrrrrrrrrrr[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:592:74  */
  assign n15878_o = ~n15877_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:52  */
  assign n15879_o = n15878_o & n15876_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:23  */
  assign n15881_o = tid[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:31  */
  assign n15882_o = tid_delay[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:604:38  */
  assign n15883_o = delay_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:601:16  */
  assign n15885_o = n15882_o ? 1'b0 : n15883_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:599:16  */
  assign n15887_o = n15881_o ? 1'b1 : n15885_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:608:28  */
  assign n15888_o = vm_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:609:44  */
  assign n15889_o = data_model_r[31:30];
  /* ../../HW/src/pcore/instr_fetch.vhd:610:34  */
  assign n15890_o = tid_rrrrrrrrrrr[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:613:30  */
  assign n15891_o = ~ready;
  /* ../../HW/src/pcore/instr_fetch.vhd:616:32  */
  assign n15892_o = pc_r[10:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:617:36  */
  assign n15893_o = busy_r[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:618:27  */
  assign n15894_o = tid[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:35  */
  assign n15895_o = tid_delay[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:623:42  */
  assign n15896_o = delay_r[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:620:20  */
  assign n15898_o = n15895_o ? 1'b0 : n15896_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:618:20  */
  assign n15900_o = n15894_o ? 1'b1 : n15898_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15901_o = n15890_o ? next_addr : n15892_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15902_o = n15890_o ? n15891_o : n15893_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:610:16  */
  assign n15904_o = n15890_o ? 1'b1 : n15900_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15905_o = n15879_o ? 1'b0 : n15853_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15906_o = n15879_o ? task_start_addr_r : n15901_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15908_o = n15879_o ? 1'b1 : n15902_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15909_o = n15879_o ? n15887_o : n15904_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15910_o = n15879_o ? task_vm_r : n15888_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15911_o = n15879_o ? task2_data_model_r : n15889_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:592:12  */
  assign n15914_o = n15879_o ? 1'b1 : 1'b0;
  assign n15915_o = iregister_auto_r[447:420];
  /* ../../HW/src/pcore/instr_fetch.vhd:633:12  */
  assign n15916_o = n15914_o ? task_iregister_auto_r : n15915_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:37  */
  assign n15917_o = ~n15909_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:26  */
  assign n15918_o = n15917_o & n15908_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:54  */
  assign n15919_o = next_tid[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:636:57  */
  assign n15920_o = ~n15919_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:42  */
  assign n15921_o = n15920_o & n15918_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:636:12  */
  assign n15924_o = n15921_o ? 1'b1 : 1'b0;
  assign n15925_o = {n14986_o, n15048_o, n15110_o, n15172_o, n15234_o, n15296_o, n15358_o, n15420_o, n15482_o, n15544_o, n15606_o, n15668_o, n15730_o, n15792_o, n15854_o, n15906_o};
  assign n15927_o = {n15908_o, n15856_o, n15794_o, n15732_o, n15670_o, n15608_o, n15546_o, n15484_o, n15422_o, n15360_o, n15298_o, n15236_o, n15174_o, n15112_o, n15050_o, n14988_o};
  assign n15929_o = {n15910_o, n15858_o, n15796_o, n15734_o, n15672_o, n15610_o, n15548_o, n15486_o, n15424_o, n15362_o, n15300_o, n15238_o, n15176_o, n15114_o, n15052_o, n14990_o};
  assign n15932_o = {n15911_o, n15859_o, n15797_o, n15735_o, n15673_o, n15611_o, n15549_o, n15487_o, n15425_o, n15363_o, n15301_o, n15239_o, n15177_o, n15115_o, n15053_o, n14991_o};
  assign n15935_o = {n15916_o, n15864_o, n15802_o, n15740_o, n15678_o, n15616_o, n15554_o, n15492_o, n15430_o, n15368_o, n15306_o, n15244_o, n15182_o, n15120_o, n15058_o, n14996_o};
  assign n15938_o = {n14989_o, n15051_o, n15113_o, n15175_o, n15237_o, n15299_o, n15361_o, n15423_o, n15485_o, n15547_o, n15609_o, n15671_o, n15733_o, n15795_o, n15857_o, n15909_o};
  assign n15940_o = {n15924_o, n15872_o, n15810_o, n15748_o, n15686_o, n15624_o, n15562_o, n15500_o, n15438_o, n15376_o, n15314_o, n15252_o, n15190_o, n15128_o, n15066_o, n15004_o};
  assign n15947_o = {n15905_o, n15848_o, n15786_o, n15724_o, n15662_o, n15600_o, n15538_o, n15476_o, n15414_o, n15352_o, n15290_o, n15228_o, n15166_o, n15104_o, n15042_o, n14980_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:652:30  */
  assign n16036_o = rom_data_in[127:48];
  /* ../../HW/src/pcore/instr_fetch.vhd:653:31  */
  assign n16037_o = rom_data_in[47:16];
  /* ../../HW/src/pcore/instr_fetch.vhd:654:32  */
  assign n16038_o = rom_data_in[15:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:662:12  */
  assign n16042_o = ~reset_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:693:51  */
  assign n16044_o = ctrl_instruction[15:11];
  /* ../../HW/src/pcore/instr_fetch.vhd:693:109  */
  assign n16046_o = n16044_o != 5'b00000;
  /* ../../HW/src/pcore/instr_fetch.vhd:693:31  */
  assign n16047_o = n16046_o & tid_valid_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:693:9  */
  assign n16050_o = n16047_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:699:42  */
  assign n16051_o = ctrl_instruction[15:11];
  /* ../../HW/src/pcore/instr_fetch.vhd:700:45  */
  assign n16052_o = ctrl_instruction[10:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:726:106  */
  assign n16053_o = instruction_addr_rr[10:1];
  /* ../../HW/src/pcore/instr_fetch.vhd:726:139  */
  assign n16055_o = n16053_o + 10'b0000000001;
  /* ../../HW/src/pcore/instr_fetch.vhd:734:9  */
  assign n16057_o = ctrl_jump ? ctrl_goto_addr_rrrrrrrr : ctrl_next_addr_rrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:732:9  */
  assign n16059_o = ctrl_ret_func ? 11'b00000000000 : n16057_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:740:32  */
  assign n16061_o = ctrl_opcode_rrrrrrrr == 5'b00001;
  /* ../../HW/src/pcore/instr_fetch.vhd:740:54  */
  assign n16062_o = got_control_rrrrrrrr & n16061_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:740:9  */
  assign n16065_o = n16062_o ? 1'b1 : 1'b0;
  assign n16080_o = {n16055_o, 1'b0};
  /* ../../HW/src/pcore/instr_fetch.vhd:758:13  */
  assign n16161_o = ctrl_opcode_rrrrrrrr == 5'b00001;
  /* ../../HW/src/pcore/instr_fetch.vhd:761:13  */
  assign n16163_o = ctrl_opcode_rrrrrrrr == 5'b00010;
  /* ../../HW/src/pcore/instr_fetch.vhd:765:42  */
  assign n16164_o = i_y_neg_in | i_y_zero_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:764:13  */
  assign n16166_o = ctrl_opcode_rrrrrrrr == 5'b00011;
  /* ../../HW/src/pcore/instr_fetch.vhd:768:31  */
  assign n16167_o = ~i_y_neg_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:768:52  */
  assign n16168_o = ~i_y_zero_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:768:47  */
  assign n16169_o = n16167_o & n16168_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:767:13  */
  assign n16171_o = ctrl_opcode_rrrrrrrr == 5'b00100;
  /* ../../HW/src/pcore/instr_fetch.vhd:771:31  */
  assign n16172_o = ~i_y_neg_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:770:13  */
  assign n16174_o = ctrl_opcode_rrrrrrrr == 5'b00101;
  /* ../../HW/src/pcore/instr_fetch.vhd:773:13  */
  assign n16176_o = ctrl_opcode_rrrrrrrr == 5'b00110;
  /* ../../HW/src/pcore/instr_fetch.vhd:777:30  */
  assign n16177_o = ~i_y_zero_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:776:13  */
  assign n16179_o = ctrl_opcode_rrrrrrrr == 5'b00111;
  /* ../../HW/src/pcore/instr_fetch.vhd:779:13  */
  assign n16181_o = ctrl_opcode_rrrrrrrr == 5'b01000;
  assign n16182_o = {n16181_o, n16179_o, n16176_o, n16174_o, n16171_o, n16166_o, n16163_o, n16161_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:757:9  */
  always @*
    case (n16182_o)
      8'b10000000: n16186_o = 1'b1;
      8'b01000000: n16186_o = n16177_o;
      8'b00100000: n16186_o = i_y_zero_in;
      8'b00010000: n16186_o = n16172_o;
      8'b00001000: n16186_o = n16169_o;
      8'b00000100: n16186_o = n16164_o;
      8'b00000010: n16186_o = i_y_neg_in;
      8'b00000001: n16186_o = 1'b0;
      default: n16186_o = 1'b0;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:757:9  */
  always @*
    case (n16182_o)
      8'b10000000: n16196_o = 1'b0;
      8'b01000000: n16196_o = 1'b0;
      8'b00100000: n16196_o = 1'b0;
      8'b00010000: n16196_o = 1'b0;
      8'b00001000: n16196_o = 1'b0;
      8'b00000100: n16196_o = 1'b0;
      8'b00000010: n16196_o = 1'b0;
      8'b00000001: n16196_o = 1'b1;
      default: n16196_o = 1'b0;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:756:5  */
  assign n16198_o = got_control_rrrrrrrr ? n16186_o : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:756:5  */
  assign n16200_o = got_control_rrrrrrrr ? n16196_o : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:795:12  */
  assign n16204_o = ~reset_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:808:12  */
  assign n16215_o = ~reset_in;
  /* ../../HW/src/pcore/instr_fetch.vhd:814:26  */
  assign n16217_o = ~task_lockstep_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16219_o = task_pcore_curr_r == 5'b00000;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16222_o = n16219_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16224_o = task_pcore_curr_r == 5'b00001;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16227_o = n16224_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16229_o = task_pcore_curr_r == 5'b00010;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16232_o = n16229_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16234_o = task_pcore_curr_r == 5'b00011;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16237_o = n16234_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16239_o = task_pcore_curr_r == 5'b00100;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16242_o = n16239_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16244_o = task_pcore_curr_r == 5'b00101;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16247_o = n16244_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16249_o = task_pcore_curr_r == 5'b00110;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16252_o = n16249_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:34  */
  assign n16254_o = task_pcore_curr_r == 5'b00111;
  /* ../../HW/src/pcore/instr_fetch.vhd:816:14  */
  assign n16257_o = n16254_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16259_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00000);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16262_o = n16259_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16264_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00001);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16267_o = n16264_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16269_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00010);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16272_o = n16269_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16274_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00011);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16277_o = n16274_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16279_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00100);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16282_o = n16279_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16284_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00101);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16287_o = n16284_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16289_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00110);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16292_o = n16289_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr_fetch.vhd:824:34  */
  assign n16294_o = $unsigned(task_pcore_max_r) >= $unsigned(5'b00111);
  /* ../../HW/src/pcore/instr_fetch.vhd:824:14  */
  assign n16297_o = n16294_o ? 1'b1 : 1'b0;
  assign n16298_o = {n16297_o, n16292_o, n16287_o, n16282_o, n16277_o, n16272_o, n16267_o, n16262_o};
  assign n16299_o = {n16257_o, n16252_o, n16247_o, n16242_o, n16237_o, n16232_o, n16227_o, n16222_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:814:8  */
  assign n16300_o = n16217_o ? n16299_o : n16298_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16308_q <= 176'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n16308_q <= n15925_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16309_q <= 16'b0000000000000000;
    else
      n16309_q <= n15927_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16310_q <= 16'b0000000000000000;
    else
      n16310_q <= n15929_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16311_q <= 16'b0000000000000000;
    else
      n16311_q <= vm_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16312_q <= 32'b00000000000000000000000000000000;
    else
      n16312_q <= n15932_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16313_q <= 32'b00000000000000000000000000000000;
    else
      n16313_q <= data_model_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16314_q <= 448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n16314_q <= n15935_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16315_q <= 448'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n16315_q <= iregister_auto_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16325_q <= 16'b0000000000000000;
    else
      n16325_q <= next_tid;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16326_q <= 1'b0;
    else
      n16326_q <= next_tid_valid;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16327_q <= 16'b0000000000000000;
    else
      n16327_q <= tid_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16328_q <= 1'b0;
    else
      n16328_q <= tid_valid_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16329_q <= 1'b0;
    else
      n16329_q <= tid_valid_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16330_q <= 16'b0000000000000000;
    else
      n16330_q <= tid_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16331_q <= 16'b0000000000000000;
    else
      n16331_q <= tid_rrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16332_q <= 16'b0000000000000000;
    else
      n16332_q <= tid_rrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16333_q <= 16'b0000000000000000;
    else
      n16333_q <= tid_rrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16334_q <= 16'b0000000000000000;
    else
      n16334_q <= tid_rrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16335_q <= 16'b0000000000000000;
    else
      n16335_q <= tid_rrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16336_q <= 16'b0000000000000000;
    else
      n16336_q <= tid_rrrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16337_q <= 16'b0000000000000000;
    else
      n16337_q <= tid_rrrrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16338_q <= 16'b0000000000000000;
    else
      n16338_q <= tid_rrrrrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16339_q <= 4'b0000;
    else
      n16339_q <= next_tid2;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16340_q <= 4'b0000;
    else
      n16340_q <= tid2_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16341_q <= 4'b0000;
    else
      n16341_q <= tid2_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16342_q <= 11'b00000000000;
    else
      n16342_q <= rom_addr;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16343_q <= 11'b00000000000;
    else
      n16343_q <= rom_addr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16344_q <= 16'b0000000000000000;
    else
      n16344_q <= n15938_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:536:5  */
  assign n16345_o = {n14332_o, n14340_o, n14348_o, n14356_o, n14364_o, n14372_o, n14380_o, n14388_o, n14396_o, n14404_o, n14412_o, n14420_o, n14428_o, n14436_o, n14444_o, n14452_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16346_q <= 2'b00;
    else
      n16346_q <= busy2;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16347_q <= 16'b0000000000000000;
    else
      n16347_q <= n15940_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16348_q <= 80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n16348_q <= mu_instruction;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16349_q <= 32'b00000000000000000000000000000000;
    else
      n16349_q <= imu_instruction;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16350_q <= 1'b0;
    else
      n16350_q <= n14676_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  always @(posedge clock_in or posedge n14668_o)
    if (n14668_o)
      n16351_q <= 1'b0;
    else
      n16351_q <= n14683_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16352_o = task_in ? task_start_addr_in : task_start_addr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16353_q <= 11'b00000000000;
    else
      n16353_q <= n16352_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16354_o = task_in ? task_pcore_max_in : task_pcore_max_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16355_q <= 5'b00000;
    else
      n16355_q <= n16354_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16356_q <= 5'b00000;
    else
      n16356_q <= n14941_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16357_o = task_in ? task_tid_mask : task_tid_mask_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16358_q <= 16'b1111111111111111;
    else
      n16358_q <= n16357_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16359_o = task_in ? task_lockstep_in : task_lockstep_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16360_q <= 1'b0;
    else
      n16360_q <= n16359_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16361_q <= 16'b0000000000000000;
    else
      n16361_q <= n15947_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16362_o = task_in ? task_vm_in : task_vm_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16363_q <= 1'b0;
    else
      n16363_q <= n16362_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16364_o = task_in ? task_iregister_auto_in : task_iregister_auto_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16365_q <= 28'b0000000000000000000000000000;
    else
      n16365_q <= n16364_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16366_o = task_in ? task_data_model_in : task2_data_model_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16367_q <= 2'b00;
    else
      n16367_q <= n16366_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:799:5  */
  always @(posedge clock_in or posedge n16204_o)
    if (n16204_o)
      n16368_q <= 11'b00000000000;
    else
      n16368_q <= rom_addr_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:799:5  */
  always @(posedge clock_in or posedge n16204_o)
    if (n16204_o)
      n16369_q <= 11'b00000000000;
    else
      n16369_q <= instruction_addr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:659:1  */
  assign n16370_o = ~n16042_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  assign n16371_o = n16370_o ? n16050_o : got_control_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in)
    n16372_q <= n16371_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16373_q <= 1'b0;
    else
      n16373_q <= got_control_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16374_q <= 1'b0;
    else
      n16374_q <= got_control_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16375_q <= 1'b0;
    else
      n16375_q <= got_control_rrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16376_q <= 1'b0;
    else
      n16376_q <= got_control_rrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16377_q <= 1'b0;
    else
      n16377_q <= got_control_rrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16378_q <= 1'b0;
    else
      n16378_q <= got_control_rrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16379_q <= 1'b0;
    else
      n16379_q <= got_control_rrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:659:1  */
  assign n16380_o = ~n16042_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  assign n16381_o = n16380_o ? n16051_o : ctrl_opcode_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in)
    n16382_q <= n16381_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:659:1  */
  assign n16383_o = ~n16042_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  assign n16384_o = n16383_o ? n16052_o : ctrl_goto_addr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in)
    n16385_q <= n16384_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16386_q <= 5'b00000;
    else
      n16386_q <= ctrl_opcode_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16387_q <= 11'b00000000000;
    else
      n16387_q <= ctrl_goto_addr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16388_q <= 5'b00000;
    else
      n16388_q <= ctrl_opcode_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16389_q <= 11'b00000000000;
    else
      n16389_q <= ctrl_goto_addr_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16390_q <= 11'b00000000000;
    else
      n16390_q <= n16080_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16391_q <= 11'b00000000000;
    else
      n16391_q <= ctrl_next_addr_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16392_q <= 11'b00000000000;
    else
      n16392_q <= ctrl_next_addr_rr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16393_q <= 11'b00000000000;
    else
      n16393_q <= ctrl_next_addr_rrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16394_q <= 11'b00000000000;
    else
      n16394_q <= ctrl_next_addr_rrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16395_q <= 11'b00000000000;
    else
      n16395_q <= n16059_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16396_q <= 1'b0;
    else
      n16396_q <= n16065_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16397_q <= 5'b00000;
    else
      n16397_q <= ctrl_opcode_rrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16398_q <= 5'b00000;
    else
      n16398_q <= ctrl_opcode_rrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16399_q <= 5'b00000;
    else
      n16399_q <= ctrl_opcode_rrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16400_q <= 5'b00000;
    else
      n16400_q <= ctrl_opcode_rrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16401_q <= 5'b00000;
    else
      n16401_q <= ctrl_opcode_rrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16402_q <= 11'b00000000000;
    else
      n16402_q <= ctrl_goto_addr_rrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16403_q <= 11'b00000000000;
    else
      n16403_q <= ctrl_goto_addr_rrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16404_q <= 11'b00000000000;
    else
      n16404_q <= ctrl_goto_addr_rrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16405_q <= 11'b00000000000;
    else
      n16405_q <= ctrl_goto_addr_rrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:692:5  */
  always @(posedge clock_in or posedge n16042_o)
    if (n16042_o)
      n16406_q <= 11'b00000000000;
    else
      n16406_q <= ctrl_goto_addr_rrrrrrr;
  /* ../../HW/src/pcore/instr_fetch.vhd:812:5  */
  always @(posedge clock_in or posedge n16215_o)
    if (n16215_o)
      n16407_q <= 8'b00000000;
    else
      n16407_q <= n16300_o;
  /* ../../HW/src/pcore/instr_fetch.vhd:812:5  */
  always @(posedge clock_in or posedge n16215_o)
    if (n16215_o)
      n16408_q <= 8'b00000000;
    else
      n16408_q <= instruction_pcore_enable_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16409_q <= 1'b0;
    else
      n16409_q <= tid_vm;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16410_q <= 1'b0;
    else
      n16410_q <= tid_vm_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16411_q <= 2'b00;
    else
      n16411_q <= task_data_model;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16412_q <= 2'b00;
    else
      n16412_q <= task_data_model_r;
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  always @(posedge clock_in or posedge n14918_o)
    if (n14918_o)
      n16413_q <= 28'b0000000000000000000000000000;
    else
      n16413_q <= tid_iregister_auto;
  /* ../../HW/src/pcore/instr_fetch.vhd:536:5  */
  assign n16414_o = {n14308_o, n14301_o};
  /* ../../HW/src/pcore/instr_fetch.vhd:513:40  */
  assign n16415_o = iregister_auto_rr[27:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:512:34  */
  assign n16416_o = iregister_auto_rr[55:28];
  /* ../../HW/src/pcore/instr_fetch.vhd:504:1  */
  assign n16417_o = iregister_auto_rr[83:56];
  /* ../../HW/src/pcore/instr_fetch.vhd:504:1  */
  assign n16418_o = iregister_auto_rr[111:84];
  /* ../../HW/src/pcore/instr_fetch.vhd:383:96  */
  assign n16419_o = iregister_auto_rr[139:112];
  /* ../../HW/src/pcore/instr_fetch.vhd:382:1  */
  assign n16420_o = iregister_auto_rr[167:140];
  /* ../../HW/src/pcore/instr_fetch.vhd:68:16  */
  assign n16421_o = iregister_auto_rr[195:168];
  /* ../../HW/src/pcore/instr_fetch.vhd:67:16  */
  assign n16422_o = iregister_auto_rr[223:196];
  /* ../../HW/src/pcore/instr_fetch.vhd:62:16  */
  assign n16423_o = iregister_auto_rr[251:224];
  /* ../../HW/src/pcore/instr_fetch.vhd:61:16  */
  assign n16424_o = iregister_auto_rr[279:252];
  /* ../../HW/src/pcore/instr_fetch.vhd:57:16  */
  assign n16425_o = iregister_auto_rr[307:280];
  /* ../../HW/src/pcore/instr_fetch.vhd:56:16  */
  assign n16426_o = iregister_auto_rr[335:308];
  /* ../../HW/src/pcore/instr_fetch.vhd:55:16  */
  assign n16427_o = iregister_auto_rr[363:336];
  /* ../../HW/src/pcore/instr_fetch.vhd:54:16  */
  assign n16428_o = iregister_auto_rr[391:364];
  /* ../../HW/src/pcore/instr_fetch.vhd:53:16  */
  assign n16429_o = iregister_auto_rr[419:392];
  /* ../../HW/src/pcore/instr_fetch.vhd:52:16  */
  assign n16430_o = iregister_auto_rr[447:420];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  assign n16431_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  always @*
    case (n16431_o)
      2'b00: n16432_o = n16415_o;
      2'b01: n16432_o = n16416_o;
      2'b10: n16432_o = n16417_o;
      2'b11: n16432_o = n16418_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  assign n16433_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  always @*
    case (n16433_o)
      2'b00: n16434_o = n16419_o;
      2'b01: n16434_o = n16420_o;
      2'b10: n16434_o = n16421_o;
      2'b11: n16434_o = n16422_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  assign n16435_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  always @*
    case (n16435_o)
      2'b00: n16436_o = n16423_o;
      2'b01: n16436_o = n16424_o;
      2'b10: n16436_o = n16425_o;
      2'b11: n16436_o = n16426_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  assign n16437_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  always @*
    case (n16437_o)
      2'b00: n16438_o = n16427_o;
      2'b01: n16438_o = n16428_o;
      2'b10: n16438_o = n16429_o;
      2'b11: n16438_o = n16430_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  assign n16439_o = tid2_r[3:2];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  always @*
    case (n16439_o)
      2'b00: n16440_o = n16432_o;
      2'b01: n16440_o = n16434_o;
      2'b10: n16440_o = n16436_o;
      2'b11: n16440_o = n16438_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:360:40  */
  assign n16441_o = vm_rr[0];
  /* ../../HW/src/pcore/instr_fetch.vhd:360:41  */
  assign n16442_o = vm_rr[1];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16443_o = vm_rr[2];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16444_o = vm_rr[3];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16445_o = vm_rr[4];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16446_o = vm_rr[5];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16447_o = vm_rr[6];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16448_o = vm_rr[7];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16449_o = vm_rr[8];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16450_o = vm_rr[9];
  /* ../../HW/src/pcore/instr_fetch.vhd:449:9  */
  assign n16451_o = vm_rr[10];
  assign n16452_o = vm_rr[11];
  /* ../../HW/src/pcore/instr_fetch.vhd:806:1  */
  assign n16453_o = vm_rr[12];
  assign n16454_o = vm_rr[13];
  /* ../../HW/src/pcore/instr_fetch.vhd:793:1  */
  assign n16455_o = vm_rr[14];
  assign n16456_o = vm_rr[15];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  assign n16457_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  always @*
    case (n16457_o)
      2'b00: n16458_o = n16441_o;
      2'b01: n16458_o = n16442_o;
      2'b10: n16458_o = n16443_o;
      2'b11: n16458_o = n16444_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  assign n16459_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  always @*
    case (n16459_o)
      2'b00: n16460_o = n16445_o;
      2'b01: n16460_o = n16446_o;
      2'b10: n16460_o = n16447_o;
      2'b11: n16460_o = n16448_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  assign n16461_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  always @*
    case (n16461_o)
      2'b00: n16462_o = n16449_o;
      2'b01: n16462_o = n16450_o;
      2'b10: n16462_o = n16451_o;
      2'b11: n16462_o = n16452_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  assign n16463_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  always @*
    case (n16463_o)
      2'b00: n16464_o = n16453_o;
      2'b01: n16464_o = n16454_o;
      2'b10: n16464_o = n16455_o;
      2'b11: n16464_o = n16456_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  assign n16465_o = tid2_r[3:2];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  always @*
    case (n16465_o)
      2'b00: n16466_o = n16458_o;
      2'b01: n16466_o = n16460_o;
      2'b10: n16466_o = n16462_o;
      2'b11: n16466_o = n16464_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:362:16  */
  assign n16467_o = data_model_rr[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:362:17  */
  assign n16468_o = data_model_rr[3:2];
  /* ../../HW/src/pcore/instr_fetch.vhd:528:1  */
  assign n16469_o = data_model_rr[5:4];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16470_o = data_model_rr[7:6];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16471_o = data_model_rr[9:8];
  /* ../../HW/src/pcore/instr_fetch.vhd:528:1  */
  assign n16472_o = data_model_rr[11:10];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16473_o = data_model_rr[13:12];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16474_o = data_model_rr[15:14];
  /* ../../HW/src/pcore/instr_fetch.vhd:528:1  */
  assign n16475_o = data_model_rr[17:16];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16476_o = data_model_rr[19:18];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16477_o = data_model_rr[21:20];
  /* ../../HW/src/pcore/instr_fetch.vhd:528:1  */
  assign n16478_o = data_model_rr[23:22];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16479_o = data_model_rr[25:24];
  /* ../../HW/src/pcore/instr_fetch.vhd:562:5  */
  assign n16480_o = data_model_rr[27:26];
  /* ../../HW/src/pcore/instr_fetch.vhd:528:1  */
  assign n16481_o = data_model_rr[29:28];
  assign n16482_o = data_model_rr[31:30];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  assign n16483_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  always @*
    case (n16483_o)
      2'b00: n16484_o = n16467_o;
      2'b01: n16484_o = n16468_o;
      2'b10: n16484_o = n16469_o;
      2'b11: n16484_o = n16470_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  assign n16485_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  always @*
    case (n16485_o)
      2'b00: n16486_o = n16471_o;
      2'b01: n16486_o = n16472_o;
      2'b10: n16486_o = n16473_o;
      2'b11: n16486_o = n16474_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  assign n16487_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  always @*
    case (n16487_o)
      2'b00: n16488_o = n16475_o;
      2'b01: n16488_o = n16476_o;
      2'b10: n16488_o = n16477_o;
      2'b11: n16488_o = n16478_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  assign n16489_o = tid2_r[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  always @*
    case (n16489_o)
      2'b00: n16490_o = n16479_o;
      2'b01: n16490_o = n16480_o;
      2'b10: n16490_o = n16481_o;
      2'b11: n16490_o = n16482_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  assign n16491_o = tid2_r[3:2];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  always @*
    case (n16491_o)
      2'b00: n16492_o = n16484_o;
      2'b01: n16492_o = n16486_o;
      2'b10: n16492_o = n16488_o;
      2'b11: n16492_o = n16490_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:364:33  */
  assign n16493_o = pc_r[10:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:364:34  */
  assign n16494_o = pc_r[21:11];
  assign n16495_o = pc_r[32:22];
  assign n16496_o = pc_r[43:33];
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n16497_o = pc_r[54:44];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n16498_o = pc_r[65:55];
  assign n16499_o = pc_r[76:66];
  assign n16500_o = pc_r[87:77];
  assign n16501_o = pc_r[98:88];
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n16502_o = pc_r[109:99];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n16503_o = pc_r[120:110];
  assign n16504_o = pc_r[131:121];
  assign n16505_o = pc_r[142:132];
  assign n16506_o = pc_r[153:143];
  /* ../../HW/src/pcore/instr_fetch.vhd:583:8  */
  assign n16507_o = pc_r[164:154];
  /* ../../HW/src/pcore/instr_fetch.vhd:571:9  */
  assign n16508_o = pc_r[175:165];
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  assign n16509_o = n14290_o[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  always @*
    case (n16509_o)
      2'b00: n16510_o = n16493_o;
      2'b01: n16510_o = n16494_o;
      2'b10: n16510_o = n16495_o;
      2'b11: n16510_o = n16496_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  assign n16511_o = n14290_o[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  always @*
    case (n16511_o)
      2'b00: n16512_o = n16497_o;
      2'b01: n16512_o = n16498_o;
      2'b10: n16512_o = n16499_o;
      2'b11: n16512_o = n16500_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  assign n16513_o = n14290_o[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  always @*
    case (n16513_o)
      2'b00: n16514_o = n16501_o;
      2'b01: n16514_o = n16502_o;
      2'b10: n16514_o = n16503_o;
      2'b11: n16514_o = n16504_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  assign n16515_o = n14290_o[1:0];
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  always @*
    case (n16515_o)
      2'b00: n16516_o = n16505_o;
      2'b01: n16516_o = n16506_o;
      2'b10: n16516_o = n16507_o;
      2'b11: n16516_o = n16508_o;
    endcase
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  assign n16517_o = n14290_o[3:2];
  /* ../../HW/src/pcore/instr_fetch.vhd:366:17  */
  always @*
    case (n16517_o)
      2'b00: n16518_o = n16510_o;
      2'b01: n16518_o = n16512_o;
      2'b10: n16518_o = n16514_o;
      2'b11: n16518_o = n16516_o;
    endcase
endmodule

module rom
  (input  clock_in,
   input  reset_in,
   input  [10:0] rdaddress_in,
   input  [10:0] rdaddress_plus_2_in,
   input  wren_in,
   input  [10:0] wraddress_in,
   input  [63:0] wrdata_in,
   output [127:0] instruction_out);
  wire [9:0] address;
  wire [127:0] q;
  wire [15:0] byteena;
  wire [9:0] n14216_o;
  wire n14217_o;
  wire n14218_o;
  wire n14219_o;
  wire n14220_o;
  wire n14221_o;
  wire n14222_o;
  wire n14223_o;
  wire n14224_o;
  wire n14225_o;
  wire n14226_o;
  wire n14227_o;
  wire n14228_o;
  wire n14229_o;
  wire n14230_o;
  wire n14231_o;
  wire n14232_o;
  wire [3:0] n14233_o;
  wire [3:0] n14234_o;
  wire [7:0] n14235_o;
  wire n14236_o;
  wire n14237_o;
  wire n14238_o;
  wire n14239_o;
  wire n14240_o;
  wire n14241_o;
  wire n14242_o;
  wire n14243_o;
  wire [3:0] n14244_o;
  wire [3:0] n14245_o;
  wire [7:0] n14246_o;
  wire [9:0] n14247_o;
  wire [9:0] n14248_o;
  wire [15:0] n14249_o;
  wire [15:0] n14251_o;
  wire [127:0] n14253_o;
  wire [127:0] ram_i_n14254;
  wire [127:0] ram_i_q_a;
  assign instruction_out = q;
  /* ../../HW/src/pcore/rom.vhd:72:8  */
  assign address = n14248_o; // (signal)
  /* ../../HW/src/pcore/rom.vhd:73:8  */
  assign q = ram_i_n14254; // (signal)
  /* ../../HW/src/pcore/rom.vhd:76:8  */
  assign byteena = n14251_o; // (signal)
  /* ../../HW/src/pcore/rom.vhd:85:28  */
  assign n14216_o = wraddress_in[10:1];
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14217_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14218_o = ~n14217_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14219_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14220_o = ~n14219_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14221_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14222_o = ~n14221_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14223_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14224_o = ~n14223_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14225_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14226_o = ~n14225_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14227_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14228_o = ~n14227_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14229_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14230_o = ~n14229_o;
  /* ../../HW/src/pcore/rom.vhd:86:86  */
  assign n14231_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:86:70  */
  assign n14232_o = ~n14231_o;
  /* ../../HW/src/dp/dp_sink.vhd:755:1  */
  assign n14233_o = {n14218_o, n14220_o, n14222_o, n14224_o};
  assign n14234_o = {n14226_o, n14228_o, n14230_o, n14232_o};
  /* ../../HW/src/dp/dp_sink.vhd:755:1  */
  assign n14235_o = {n14233_o, n14234_o};
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14236_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14237_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14238_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14239_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14240_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14241_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14242_o = wraddress_in[0];
  /* ../../HW/src/pcore/rom.vhd:87:68  */
  assign n14243_o = wraddress_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14244_o = {n14236_o, n14237_o, n14238_o, n14239_o};
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14245_o = {n14240_o, n14241_o, n14242_o, n14243_o};
  /* ../../HW/src/dp/dp_sink.vhd:426:1  */
  assign n14246_o = {n14244_o, n14245_o};
  /* ../../HW/src/pcore/rom.vhd:89:28  */
  assign n14247_o = rdaddress_in[10:1];
  /* ../../HW/src/pcore/rom.vhd:84:1  */
  assign n14248_o = wren_in ? n14216_o : n14247_o;
  /* ../../HW/src/dp/dp_sink.vhd:426:1  */
  assign n14249_o = {n14235_o, n14246_o};
  /* ../../HW/src/pcore/rom.vhd:84:1  */
  assign n14251_o = wren_in ? n14249_o : 16'b0000000000000000;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14253_o = {wrdata_in, wrdata_in};
  /* ../../HW/src/pcore/rom.vhd:111:13  */
  assign ram_i_n14254 = ram_i_q_a; // (signal)
  /* ../../HW/src/pcore/rom.vhd:98:1  */
  spram_be_1024_10_128 ram_i (
    .address_a(address),
    .clock0(clock_in),
    .data_a(n14253_o),
    .wren_a(wren_in),
    .byteena_a(byteena),
    .q_a(ram_i_q_a));
endmodule

module adder_12
  (input  [11:0] x_in,
   input  [11:0] y_in,
   input  add_sub_in,
   output [11:0] z_out);
  wire [11:0] x;
  wire [11:0] y;
  wire [11:0] z;
  wire [11:0] n14209_o;
  wire [11:0] n14210_o;
  wire [11:0] n14211_o;
  assign z_out = z;
  /* ../../HW/src/util/adder.vhd:38:8  */
  assign x = x_in; // (signal)
  /* ../../HW/src/util/adder.vhd:39:8  */
  assign y = y_in; // (signal)
  /* ../../HW/src/util/adder.vhd:40:8  */
  assign z = n14211_o; // (signal)
  /* ../../HW/src/util/adder.vhd:52:14  */
  assign n14209_o = x + y;
  /* ../../HW/src/util/adder.vhd:54:14  */
  assign n14210_o = x - y;
  /* ../../HW/src/util/adder.vhd:51:4  */
  assign n14211_o = add_sub_in ? n14209_o : n14210_o;
endmodule

module multiplier_12_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clock_in,
   input  reset_in,
   input  [11:0] x_in,
   input  [11:0] y_in,
   output [23:0] z_out);
  wire [11:0] x;
  wire [11:0] y;
  wire [23:0] z;
  wire [23:0] n14193_o;
  wire [23:0] n14194_o;
  wire [23:0] n14195_o;
  assign z_out = z;
  /* ../../HW/src/util/multiplier.vhd:43:8  */
  assign x = x_in; // (signal)
  /* ../../HW/src/util/multiplier.vhd:44:8  */
  assign y = y_in; // (signal)
  /* ../../HW/src/util/multiplier.vhd:45:8  */
  assign z = n14195_o; // (signal)
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n14193_o = {{12{x[11]}}, x}; // sext
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n14194_o = {{12{y[11]}}, y}; // sext
  /* ../../HW/src/util/multiplier.vhd:51:7  */
  assign n14195_o = n14193_o * n14194_o; // smul
endmodule

module spram_512_9_24
  (input  [8:0] address_a,
   input  clock0,
   input  [23:0] data_a,
   input  wren_a,
   output [23:0] q_a);
  wire [8:0] address_r;
  reg [8:0] n14189_q;
  wire [23:0] n14190_data; // mem_rd
  assign q_a = n14190_data;
  /* ../../HW/platform/simulation/SPRAM.vhd:50:8  */
  assign address_r = n14189_q; // (signal)
  /* ../../HW/platform/simulation/SPRAM.vhd:56:7  */
  always @(posedge clock0)
    n14189_q <= address_a;
  /* ../../HW/platform/simulation/SPRAM.vhd:41:8  */
  reg [23:0] ram[511:0] ; // memory
  assign n14190_data = ram[address_r];
  always @(posedge clock0)
    if (wren_a)
      ram[address_a] <= data_a;
  /* ../../HW/platform/simulation/SPRAM.vhd:65:15  */
  /* ../../HW/platform/simulation/SPRAM.vhd:58:17  */
endmodule

module dp_sink_3_32_1_9_40623dc9948b5e96ae4a8c3b66bafc8116c42db3
  (input  clock_in,
   input  reset_in,
   input  bus_wait_request_in,
   input  [2:0] wr_req_in,
   input  [2:0] wr_req_pending_p0_in,
   input  [2:0] wr_req_pending_p1_in,
   input  [5:0] wr_data_flow_in,
   input  [8:0] wr_vector_in,
   input  [2:0] wr_stream_in,
   input  [5:0] wr_stream_id_in,
   input  [5:0] wr_scatter_in,
   input  [11:0] wr_end_in,
   input  [95:0] wr_addr_in,
   input  [2:0] wr_fork_in,
   input  [2:0] wr_addr_mode_in,
   input  [2:0] wr_src_vm_in,
   input  [2:0] wr_datavalid_in,
   input  [191:0] wr_data_in,
   input  [2:0] wr_readdatavalid_in,
   input  [2:0] wr_readdatavalid_vm_in,
   input  [191:0] wr_readdata_in,
   input  [14:0] wr_burstlen_in,
   input  [5:0] wr_bus_id_in,
   input  [2:0] wr_thread_in,
   input  [5:0] wr_data_type_in,
   input  [5:0] wr_data_model_in,
   input  [17:0] wr_mcast_in,
   output [31:0] bus_addr_out,
   output bus_fork_out,
   output bus_addr_mode_out,
   output bus_vm_out,
   output [1:0] bus_data_flow_out,
   output [2:0] bus_vector_out,
   output bus_stream_out,
   output [1:0] bus_stream_id_out,
   output [1:0] bus_scatter_out,
   output [3:0] bus_end_out,
   output [5:0] bus_mcast_out,
   output bus_cs_out,
   output bus_write_out,
   output [63:0] bus_writedata_out,
   output [4:0] bus_burstlen_out,
   output [8:0] bus_burstlen2_out,
   output [4:0] bus_burstlen3_out,
   output [1:0] bus_id_out,
   output [1:0] bus_data_type_out,
   output [1:0] bus_data_model_out,
   output bus_thread_out,
   output [4:0] wr_maxburstlen_out,
   output wr_full_out,
   output [2:0] read_pending_p0_out,
   output [2:0] read_pending_p1_out);
  wire rdreq;
  wire rdreq2;
  wire empty;
  wire emptyn;
  wire empty2;
  wire [63:0] q2;
  wire [131:0] q;
  wire [131:0] q_r;
  wire valid;
  wire valid_r;
  wire valid_rr;
  wire [1:0] bus_data_flow_r;
  wire [3:0] bus_end_r;
  wire [2:0] bus_vector_r;
  wire bus_stream_r;
  wire [1:0] bus_stream_id_r;
  wire [1:0] bus_scatter_r;
  wire [31:0] bus_addr_r;
  wire bus_fork_r;
  wire bus_addr_mode_r;
  wire bus_vm_r;
  wire [63:0] bus_writedata_r;
  wire [4:0] bus_burstlen_r;
  wire [8:0] bus_burstlen2_r;
  wire [4:0] bus_burstlen3_r;
  wire [1:0] bus_id_r;
  wire bus_thread_r;
  wire [1:0] bus_data_type_r;
  wire [1:0] bus_data_model_r;
  reg [5:0] bus_mcast_r;
  wire [8:0] req_p0_0_r;
  wire [8:0] req_p0_1_r;
  wire [8:0] req_p0_2_r;
  wire [8:0] rsp_p0_0_r;
  wire [8:0] rsp_p0_1_r;
  wire [8:0] rsp_p0_2_r;
  wire [8:0] req_p1_0_r;
  wire [8:0] req_p1_1_r;
  wire [8:0] req_p1_2_r;
  wire [8:0] rsp_p1_0_r;
  wire [8:0] rsp_p1_1_r;
  wire [8:0] rsp_p1_2_r;
  wire [8:0] usedw;
  wire [8:0] usedw2;
  wire [131:0] fifo_data;
  wire [31:0] wr_addr;
  wire wr_fork;
  wire wr_addr_mode;
  wire wr_vm;
  wire [1:0] wr_data_flow;
  wire [2:0] wr_vector;
  wire wr_stream;
  wire [1:0] wr_stream_id;
  wire [1:0] wr_scatter;
  wire [3:0] wr_end;
  wire wr_datavalid;
  wire [63:0] wr_data;
  wire [63:0] wr_data2;
  wire [4:0] wr_burstlen;
  wire [1:0] wr_bus_id;
  wire wr_thread;
  wire [1:0] wr_data_type;
  wire [1:0] wr_data_model;
  wire [5:0] wr_mcast;
  wire wr_req;
  wire [2:0] wr_req2;
  wire wr_req2_all;
  wire [2:0] read_pending_p0_r;
  wire [2:0] read_pending_p1_r;
  wire wr_full_r;
  wire [4:0] wr_maxburstlen_r;
  wire [131:0] dp_sink_fifo_i_n13300;
  wire [8:0] dp_sink_fifo_i_n13302;
  wire dp_sink_fifo_i_n13303;
  wire [131:0] dp_sink_fifo_i_q_out;
  wire [8:0] dp_sink_fifo_i_ravail_out;
  wire [8:0] dp_sink_fifo_i_wused_out;
  wire dp_sink_fifo_i_empty_out;
  wire dp_sink_fifo_i_full_out;
  wire dp_sink_fifo_i_almost_full_out;
  wire [63:0] dp_sink_fifo_i2_n13316;
  wire [8:0] dp_sink_fifo_i2_n13318;
  wire dp_sink_fifo_i2_n13319;
  wire [63:0] dp_sink_fifo_i2_q_out;
  wire [8:0] dp_sink_fifo_i2_ravail_out;
  wire [8:0] dp_sink_fifo_i2_wused_out;
  wire dp_sink_fifo_i2_empty_out;
  wire dp_sink_fifo_i2_full_out;
  wire dp_sink_fifo_i2_almost_full_out;
  wire n13332_o;
  wire n13333_o;
  wire n13334_o;
  wire n13335_o;
  wire n13336_o;
  wire n13338_o;
  wire n13339_o;
  wire n13340_o;
  wire n13341_o;
  wire n13342_o;
  wire n13343_o;
  wire n13346_o;
  wire n13347_o;
  wire n13348_o;
  wire n13349_o;
  wire n13350_o;
  wire n13351_o;
  wire n13354_o;
  wire n13355_o;
  wire n13356_o;
  wire n13357_o;
  wire n13358_o;
  wire n13359_o;
  wire n13361_o;
  wire n13362_o;
  wire n13363_o;
  wire n13364_o;
  wire n13365_o;
  wire [2:0] n13366_o;
  wire [2:0] n13367_o;
  wire n13370_o;
  wire [63:0] n13371_o;
  wire n13372_o;
  wire [63:0] n13373_o;
  wire [63:0] n13374_o;
  wire [63:0] n13375_o;
  wire [63:0] n13376_o;
  wire n13380_o;
  wire n13381_o;
  wire [63:0] n13382_o;
  wire [31:0] n13383_o;
  wire n13384_o;
  wire n13385_o;
  wire n13386_o;
  wire [1:0] n13387_o;
  wire [2:0] n13388_o;
  wire n13389_o;
  wire [1:0] n13390_o;
  wire [1:0] n13391_o;
  wire [3:0] n13392_o;
  wire [4:0] n13393_o;
  wire [1:0] n13394_o;
  wire n13395_o;
  wire [1:0] n13396_o;
  wire [1:0] n13397_o;
  wire [5:0] n13398_o;
  wire n13399_o;
  wire n13400_o;
  wire [63:0] n13401_o;
  wire [31:0] n13402_o;
  wire n13403_o;
  wire n13404_o;
  wire n13405_o;
  wire [1:0] n13406_o;
  wire [2:0] n13407_o;
  wire n13408_o;
  wire [1:0] n13409_o;
  wire [1:0] n13410_o;
  wire [3:0] n13411_o;
  wire [4:0] n13412_o;
  wire [1:0] n13413_o;
  wire n13414_o;
  wire [1:0] n13415_o;
  wire [1:0] n13416_o;
  wire [5:0] n13417_o;
  wire n13418_o;
  wire [63:0] n13419_o;
  wire [31:0] n13420_o;
  wire n13421_o;
  wire n13422_o;
  wire n13423_o;
  wire [1:0] n13424_o;
  wire [2:0] n13425_o;
  wire n13426_o;
  wire [1:0] n13427_o;
  wire [1:0] n13428_o;
  wire [3:0] n13429_o;
  wire [4:0] n13430_o;
  wire [1:0] n13431_o;
  wire n13432_o;
  wire [1:0] n13433_o;
  wire [1:0] n13434_o;
  wire [5:0] n13435_o;
  wire [31:0] n13436_o;
  wire n13437_o;
  wire n13438_o;
  wire n13439_o;
  wire [1:0] n13440_o;
  wire [2:0] n13441_o;
  wire n13442_o;
  wire [1:0] n13443_o;
  wire [1:0] n13444_o;
  wire [3:0] n13445_o;
  wire n13446_o;
  wire [63:0] n13447_o;
  wire [4:0] n13448_o;
  wire [1:0] n13449_o;
  wire n13450_o;
  wire [1:0] n13451_o;
  wire [1:0] n13452_o;
  wire [5:0] n13453_o;
  wire [31:0] n13454_o;
  wire n13455_o;
  wire n13456_o;
  wire n13457_o;
  wire [1:0] n13458_o;
  wire [2:0] n13459_o;
  wire n13460_o;
  wire [1:0] n13461_o;
  wire [1:0] n13462_o;
  wire [3:0] n13463_o;
  wire n13464_o;
  wire [63:0] n13465_o;
  wire [4:0] n13466_o;
  wire [1:0] n13467_o;
  wire n13468_o;
  wire [1:0] n13469_o;
  wire [1:0] n13470_o;
  wire [5:0] n13471_o;
  wire n13513_o;
  wire n13516_o;
  wire n13517_o;
  wire n13518_o;
  wire n13519_o;
  wire n13520_o;
  wire [8:0] n13522_o;
  wire [8:0] n13523_o;
  wire n13524_o;
  wire n13525_o;
  wire n13526_o;
  wire n13527_o;
  wire n13528_o;
  wire [8:0] n13530_o;
  wire [8:0] n13531_o;
  wire n13532_o;
  wire n13533_o;
  wire n13534_o;
  wire n13535_o;
  wire n13536_o;
  wire [8:0] n13538_o;
  wire [8:0] n13539_o;
  wire n13540_o;
  wire n13541_o;
  wire n13542_o;
  wire n13543_o;
  wire [8:0] n13545_o;
  wire [8:0] n13546_o;
  wire n13547_o;
  wire n13548_o;
  wire n13549_o;
  wire n13550_o;
  wire [8:0] n13552_o;
  wire [8:0] n13553_o;
  wire n13554_o;
  wire n13555_o;
  wire n13556_o;
  wire n13557_o;
  wire [8:0] n13559_o;
  wire [8:0] n13560_o;
  wire n13561_o;
  wire n13562_o;
  wire n13563_o;
  wire n13564_o;
  wire [8:0] n13566_o;
  wire [8:0] n13567_o;
  wire n13568_o;
  wire n13569_o;
  wire n13570_o;
  wire n13571_o;
  wire [8:0] n13573_o;
  wire [8:0] n13574_o;
  wire n13575_o;
  wire n13576_o;
  wire n13577_o;
  wire n13578_o;
  wire [8:0] n13580_o;
  wire [8:0] n13581_o;
  wire n13582_o;
  wire n13583_o;
  wire n13584_o;
  wire [8:0] n13586_o;
  wire [8:0] n13587_o;
  wire n13588_o;
  wire n13589_o;
  wire n13590_o;
  wire [8:0] n13592_o;
  wire [8:0] n13593_o;
  wire n13594_o;
  wire n13595_o;
  wire n13596_o;
  wire [8:0] n13598_o;
  wire [8:0] n13599_o;
  wire n13600_o;
  wire n13603_o;
  wire n13604_o;
  wire n13607_o;
  wire n13608_o;
  wire n13611_o;
  wire n13612_o;
  wire n13615_o;
  wire n13616_o;
  wire n13619_o;
  wire n13620_o;
  wire n13623_o;
  wire n13624_o;
  wire n13625_o;
  wire n13626_o;
  wire n13627_o;
  wire [63:0] n13628_o;
  wire [63:0] n13629_o;
  wire [31:0] n13630_o;
  wire n13631_o;
  wire n13632_o;
  wire n13633_o;
  wire [4:0] n13634_o;
  wire n13635_o;
  wire [8:0] n13637_o;
  wire [8:0] n13639_o;
  wire [8:0] n13640_o;
  wire [8:0] n13642_o;
  wire n13643_o;
  wire [4:0] n13644_o;
  wire [4:0] n13645_o;
  wire [1:0] n13646_o;
  wire n13647_o;
  wire [1:0] n13648_o;
  wire [1:0] n13649_o;
  wire [5:0] n13650_o;
  wire [2:0] n13651_o;
  wire n13652_o;
  wire [1:0] n13653_o;
  wire [1:0] n13654_o;
  wire [1:0] n13655_o;
  wire [3:0] n13656_o;
  wire [8:0] n13657_o;
  wire n13659_o;
  wire n13661_o;
  wire [8:0] n13663_o;
  wire [4:0] n13664_o;
  wire [8:0] n13666_o;
  wire n13668_o;
  wire n13670_o;
  wire [8:0] n13672_o;
  wire [4:0] n13673_o;
  wire [8:0] n13675_o;
  wire n13677_o;
  wire n13679_o;
  wire [8:0] n13681_o;
  wire [4:0] n13682_o;
  wire [8:0] n13684_o;
  wire n13686_o;
  wire [8:0] n13688_o;
  wire [4:0] n13689_o;
  wire [8:0] n13690_o;
  wire [4:0] n13691_o;
  wire [8:0] n13693_o;
  wire [4:0] n13694_o;
  wire [8:0] n13696_o;
  wire [4:0] n13697_o;
  wire [2:0] n13777_o;
  wire [2:0] n13779_o;
  wire n14050_o;
  wire [8:0] n14052_o;
  wire n14054_o;
  wire n14057_o;
  wire n14072_o;
  wire n14073_o;
  wire n14074_o;
  wire n14075_o;
  wire n14076_o;
  wire n14077_o;
  wire n14078_o;
  wire n14082_o;
  wire n14084_o;
  wire n14086_o;
  wire n14089_o;
  wire n14091_o;
  wire n14093_o;
  wire n14094_o;
  wire n14095_o;
  wire n14097_o;
  wire n14099_o;
  wire n14102_o;
  wire n14103_o;
  wire n14104_o;
  wire n14105_o;
  wire [131:0] n14109_o;
  reg [131:0] n14110_q;
  wire n14111_o;
  reg n14112_q;
  wire n14113_o;
  reg n14114_q;
  wire [1:0] n14115_o;
  reg [1:0] n14116_q;
  wire [3:0] n14117_o;
  reg [3:0] n14118_q;
  wire [2:0] n14119_o;
  reg [2:0] n14120_q;
  wire n14121_o;
  reg n14122_q;
  wire [1:0] n14123_o;
  reg [1:0] n14124_q;
  wire [1:0] n14125_o;
  reg [1:0] n14126_q;
  wire [31:0] n14127_o;
  reg [31:0] n14128_q;
  wire n14129_o;
  reg n14130_q;
  wire n14131_o;
  reg n14132_q;
  wire n14133_o;
  reg n14134_q;
  wire [63:0] n14135_o;
  reg [63:0] n14136_q;
  wire [4:0] n14137_o;
  reg [4:0] n14138_q;
  wire [8:0] n14139_o;
  reg [8:0] n14140_q;
  wire [4:0] n14141_o;
  reg [4:0] n14142_q;
  wire [1:0] n14143_o;
  reg [1:0] n14144_q;
  wire n14145_o;
  reg n14146_q;
  wire [1:0] n14147_o;
  reg [1:0] n14148_q;
  wire [1:0] n14149_o;
  reg [1:0] n14150_q;
  wire [5:0] n14151_o;
  reg [5:0] n14152_q;
  reg [8:0] n14153_q;
  reg [8:0] n14154_q;
  reg [8:0] n14155_q;
  reg [8:0] n14156_q;
  reg [8:0] n14157_q;
  reg [8:0] n14158_q;
  reg [8:0] n14159_q;
  reg [8:0] n14160_q;
  reg [8:0] n14161_q;
  reg [8:0] n14162_q;
  reg [8:0] n14163_q;
  reg [8:0] n14164_q;
  wire [131:0] n14165_o;
  wire [2:0] n14166_o;
  reg [2:0] n14167_q;
  reg [2:0] n14168_q;
  reg n14169_q;
  reg [4:0] n14170_q;
  assign bus_addr_out = bus_addr_r;
  assign bus_fork_out = bus_fork_r;
  assign bus_addr_mode_out = bus_addr_mode_r;
  assign bus_vm_out = bus_vm_r;
  assign bus_data_flow_out = bus_data_flow_r;
  assign bus_vector_out = bus_vector_r;
  assign bus_stream_out = bus_stream_r;
  assign bus_stream_id_out = bus_stream_id_r;
  assign bus_scatter_out = bus_scatter_r;
  assign bus_end_out = bus_end_r;
  assign bus_mcast_out = bus_mcast_r;
  assign bus_cs_out = valid_rr;
  assign bus_write_out = valid_rr;
  assign bus_writedata_out = bus_writedata_r;
  assign bus_burstlen_out = bus_burstlen_r;
  assign bus_burstlen2_out = bus_burstlen2_r;
  assign bus_burstlen3_out = bus_burstlen3_r;
  assign bus_id_out = bus_id_r;
  assign bus_data_type_out = bus_data_type_r;
  assign bus_data_model_out = bus_data_model_r;
  assign bus_thread_out = bus_thread_r;
  assign wr_maxburstlen_out = wr_maxburstlen_r;
  assign wr_full_out = wr_full_r;
  assign read_pending_p0_out = n13366_o;
  assign read_pending_p1_out = n13367_o;
  /* ../../HW/src/dp/dp_sink.vhd:104:8  */
  assign rdreq = n14103_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:105:8  */
  assign rdreq2 = n14104_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:107:8  */
  assign empty = dp_sink_fifo_i_n13303; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:108:8  */
  assign emptyn = n14078_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:109:8  */
  assign empty2 = dp_sink_fifo_i2_n13319; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:110:8  */
  assign q2 = dp_sink_fifo_i2_n13316; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:113:8  */
  assign q = dp_sink_fifo_i_n13300; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:114:8  */
  assign q_r = n14110_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:115:8  */
  assign valid = n14105_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:116:8  */
  assign valid_r = n14112_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:117:8  */
  assign valid_rr = n14114_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:118:8  */
  assign bus_data_flow_r = n14116_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:119:8  */
  assign bus_end_r = n14118_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:120:8  */
  assign bus_vector_r = n14120_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:121:8  */
  assign bus_stream_r = n14122_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:122:8  */
  assign bus_stream_id_r = n14124_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:123:8  */
  assign bus_scatter_r = n14126_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:124:8  */
  assign bus_addr_r = n14128_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:125:8  */
  assign bus_fork_r = n14130_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:126:8  */
  assign bus_addr_mode_r = n14132_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:127:8  */
  assign bus_vm_r = n14134_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:128:8  */
  assign bus_writedata_r = n14136_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:129:8  */
  assign bus_burstlen_r = n14138_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:130:8  */
  assign bus_burstlen2_r = n14140_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:131:8  */
  assign bus_burstlen3_r = n14142_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:132:8  */
  assign bus_id_r = n14144_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:133:8  */
  assign bus_thread_r = n14146_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:134:8  */
  assign bus_data_type_r = n14148_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:135:8  */
  assign bus_data_model_r = n14150_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:136:8  */
  always @*
    bus_mcast_r = n14152_q; // (isignal)
  initial
    bus_mcast_r = 6'b111111;
  /* ../../HW/src/dp/dp_sink.vhd:137:8  */
  assign req_p0_0_r = n14153_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:138:8  */
  assign req_p0_1_r = n14154_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:139:8  */
  assign req_p0_2_r = n14155_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:140:8  */
  assign rsp_p0_0_r = n14156_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:141:8  */
  assign rsp_p0_1_r = n14157_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:142:8  */
  assign rsp_p0_2_r = n14158_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:144:8  */
  assign req_p1_0_r = n14159_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:145:8  */
  assign req_p1_1_r = n14160_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:146:8  */
  assign req_p1_2_r = n14161_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:147:8  */
  assign rsp_p1_0_r = n14162_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:148:8  */
  assign rsp_p1_1_r = n14163_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:149:8  */
  assign rsp_p1_2_r = n14164_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:155:8  */
  assign usedw = dp_sink_fifo_i_n13302; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:156:8  */
  assign usedw2 = dp_sink_fifo_i2_n13318; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:157:8  */
  assign fifo_data = n14165_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:159:8  */
  assign wr_addr = n13454_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:160:8  */
  assign wr_fork = n13455_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:161:8  */
  assign wr_addr_mode = n13456_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:162:8  */
  assign wr_vm = n13457_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:163:8  */
  assign wr_data_flow = n13458_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:164:8  */
  assign wr_vector = n13459_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:165:8  */
  assign wr_stream = n13460_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:166:8  */
  assign wr_stream_id = n13461_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:167:8  */
  assign wr_scatter = n13462_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:168:8  */
  assign wr_end = n13463_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:169:8  */
  assign wr_datavalid = n13464_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:170:8  */
  assign wr_data = n13465_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:171:8  */
  assign wr_data2 = n13376_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:172:8  */
  assign wr_burstlen = n13466_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:173:8  */
  assign wr_bus_id = n13467_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:174:8  */
  assign wr_thread = n13468_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:175:8  */
  assign wr_data_type = n13469_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:176:8  */
  assign wr_data_model = n13470_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:177:8  */
  assign wr_mcast = n13471_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:178:8  */
  assign wr_req = n13336_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:179:8  */
  assign wr_req2 = n14166_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:180:8  */
  assign wr_req2_all = n13365_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:185:8  */
  assign read_pending_p0_r = n14167_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:186:8  */
  assign read_pending_p1_r = n14168_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:188:8  */
  assign wr_full_r = n14169_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:189:8  */
  assign wr_maxburstlen_r = n14170_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:222:16  */
  assign dp_sink_fifo_i_n13300 = dp_sink_fifo_i_q_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:224:20  */
  assign dp_sink_fifo_i_n13302 = dp_sink_fifo_i_wused_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:225:20  */
  assign dp_sink_fifo_i_n13303 = dp_sink_fifo_i_empty_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:208:1  */
  scfifo_132_9_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 dp_sink_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(fifo_data),
    .write_in(wr_req),
    .read_in(rdreq),
    .q_out(dp_sink_fifo_i_q_out),
    .ravail_out(),
    .wused_out(dp_sink_fifo_i_wused_out),
    .empty_out(dp_sink_fifo_i_empty_out),
    .full_out(),
    .almost_full_out());
  /* ../../HW/src/dp/dp_sink.vhd:244:16  */
  assign dp_sink_fifo_i2_n13316 = dp_sink_fifo_i2_q_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:246:20  */
  assign dp_sink_fifo_i2_n13318 = dp_sink_fifo_i2_wused_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:247:20  */
  assign dp_sink_fifo_i2_n13319 = dp_sink_fifo_i2_empty_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:230:1  */
  scfifo_64_9_1_5ba93c9db0cff93f52b521d7420e43f6eda2784f dp_sink_fifo_i2 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(wr_data2),
    .write_in(wr_req2_all),
    .read_in(rdreq2),
    .q_out(dp_sink_fifo_i2_q_out),
    .ravail_out(),
    .wused_out(dp_sink_fifo_i2_wused_out),
    .empty_out(dp_sink_fifo_i2_empty_out),
    .full_out(),
    .almost_full_out());
  /* ../../HW/src/dp/dp_sink.vhd:282:20  */
  assign n13332_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:282:36  */
  assign n13333_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:282:24  */
  assign n13334_o = n13332_o | n13333_o;
  /* ../../HW/src/dp/dp_sink.vhd:282:52  */
  assign n13335_o = wr_req_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:282:40  */
  assign n13336_o = n13334_o | n13335_o;
  /* ../../HW/src/dp/dp_sink.vhd:284:44  */
  assign n13338_o = wr_readdatavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:284:68  */
  assign n13339_o = req_p0_0_r != rsp_p0_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:284:96  */
  assign n13340_o = req_p1_0_r != rsp_p1_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:284:82  */
  assign n13341_o = n13339_o | n13340_o;
  /* ../../HW/src/dp/dp_sink.vhd:284:52  */
  assign n13342_o = n13341_o & n13338_o;
  /* ../../HW/src/dp/dp_sink.vhd:284:19  */
  assign n13343_o = n13342_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:286:44  */
  assign n13346_o = wr_readdatavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:286:68  */
  assign n13347_o = req_p0_1_r != rsp_p0_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:286:96  */
  assign n13348_o = req_p1_1_r != rsp_p1_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:286:82  */
  assign n13349_o = n13347_o | n13348_o;
  /* ../../HW/src/dp/dp_sink.vhd:286:52  */
  assign n13350_o = n13349_o & n13346_o;
  /* ../../HW/src/dp/dp_sink.vhd:286:19  */
  assign n13351_o = n13350_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:288:44  */
  assign n13354_o = wr_readdatavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:288:68  */
  assign n13355_o = req_p0_2_r != rsp_p0_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:288:96  */
  assign n13356_o = req_p1_2_r != rsp_p1_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:288:82  */
  assign n13357_o = n13355_o | n13356_o;
  /* ../../HW/src/dp/dp_sink.vhd:288:52  */
  assign n13358_o = n13357_o & n13354_o;
  /* ../../HW/src/dp/dp_sink.vhd:288:19  */
  assign n13359_o = n13358_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:290:23  */
  assign n13361_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:290:37  */
  assign n13362_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:290:27  */
  assign n13363_o = n13361_o | n13362_o;
  /* ../../HW/src/dp/dp_sink.vhd:290:51  */
  assign n13364_o = wr_req2[2];
  /* ../../HW/src/dp/dp_sink.vhd:290:41  */
  assign n13365_o = n13363_o | n13364_o;
  /* ../../HW/src/dp/dp_sink.vhd:292:42  */
  assign n13366_o = read_pending_p0_r | wr_req_pending_p0_in;
  /* ../../HW/src/dp/dp_sink.vhd:294:42  */
  assign n13367_o = read_pending_p1_r | wr_req_pending_p1_in;
  /* ../../HW/src/dp/dp_sink.vhd:299:14  */
  assign n13370_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:300:88  */
  assign n13371_o = wr_readdata_in[63:0];
  /* ../../HW/src/dp/dp_sink.vhd:301:17  */
  assign n13372_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:302:88  */
  assign n13373_o = wr_readdata_in[127:64];
  /* ../../HW/src/dp/dp_sink.vhd:304:88  */
  assign n13374_o = wr_readdata_in[191:128];
  /* ../../HW/src/dp/dp_sink.vhd:301:4  */
  assign n13375_o = n13372_o ? n13373_o : n13374_o;
  /* ../../HW/src/dp/dp_sink.vhd:299:4  */
  assign n13376_o = n13370_o ? n13371_o : n13375_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:13  */
  assign n13380_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:313:36  */
  assign n13381_o = wr_datavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:314:26  */
  assign n13382_o = wr_data_in[63:0];
  /* ../../HW/src/dp/dp_sink.vhd:315:26  */
  assign n13383_o = wr_addr_in[31:0];
  /* ../../HW/src/dp/dp_sink.vhd:316:26  */
  assign n13384_o = wr_src_vm_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:317:29  */
  assign n13385_o = wr_fork_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:318:36  */
  assign n13386_o = wr_addr_mode_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:319:36  */
  assign n13387_o = wr_data_flow_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:320:30  */
  assign n13388_o = wr_vector_in[2:0];
  /* ../../HW/src/dp/dp_sink.vhd:321:30  */
  assign n13389_o = wr_stream_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:322:36  */
  assign n13390_o = wr_stream_id_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:323:32  */
  assign n13391_o = wr_scatter_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:324:24  */
  assign n13392_o = wr_end_in[3:0];
  /* ../../HW/src/dp/dp_sink.vhd:325:34  */
  assign n13393_o = wr_burstlen_in[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:326:30  */
  assign n13394_o = wr_bus_id_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:327:30  */
  assign n13395_o = wr_thread_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:328:36  */
  assign n13396_o = wr_data_type_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:329:38  */
  assign n13397_o = wr_data_model_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:330:28  */
  assign n13398_o = wr_mcast_in[5:0];
  /* ../../HW/src/dp/dp_sink.vhd:331:16  */
  assign n13399_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:332:36  */
  assign n13400_o = wr_datavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:333:26  */
  assign n13401_o = wr_data_in[127:64];
  /* ../../HW/src/dp/dp_sink.vhd:334:26  */
  assign n13402_o = wr_addr_in[63:32];
  /* ../../HW/src/dp/dp_sink.vhd:335:26  */
  assign n13403_o = wr_src_vm_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:336:29  */
  assign n13404_o = wr_fork_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:337:36  */
  assign n13405_o = wr_addr_mode_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:338:36  */
  assign n13406_o = wr_data_flow_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:339:30  */
  assign n13407_o = wr_vector_in[5:3];
  /* ../../HW/src/dp/dp_sink.vhd:340:30  */
  assign n13408_o = wr_stream_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:341:36  */
  assign n13409_o = wr_stream_id_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:342:32  */
  assign n13410_o = wr_scatter_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:343:24  */
  assign n13411_o = wr_end_in[7:4];
  /* ../../HW/src/dp/dp_sink.vhd:344:34  */
  assign n13412_o = wr_burstlen_in[9:5];
  /* ../../HW/src/dp/dp_sink.vhd:345:30  */
  assign n13413_o = wr_bus_id_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:346:30  */
  assign n13414_o = wr_thread_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:347:36  */
  assign n13415_o = wr_data_type_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:348:38  */
  assign n13416_o = wr_data_model_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:349:28  */
  assign n13417_o = wr_mcast_in[11:6];
  /* ../../HW/src/dp/dp_sink.vhd:351:36  */
  assign n13418_o = wr_datavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:352:26  */
  assign n13419_o = wr_data_in[191:128];
  /* ../../HW/src/dp/dp_sink.vhd:353:26  */
  assign n13420_o = wr_addr_in[95:64];
  /* ../../HW/src/dp/dp_sink.vhd:354:26  */
  assign n13421_o = wr_src_vm_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:355:29  */
  assign n13422_o = wr_fork_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:356:36  */
  assign n13423_o = wr_addr_mode_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:357:36  */
  assign n13424_o = wr_data_flow_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:358:30  */
  assign n13425_o = wr_vector_in[8:6];
  /* ../../HW/src/dp/dp_sink.vhd:359:30  */
  assign n13426_o = wr_stream_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:360:36  */
  assign n13427_o = wr_stream_id_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:361:32  */
  assign n13428_o = wr_scatter_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:362:24  */
  assign n13429_o = wr_end_in[11:8];
  /* ../../HW/src/dp/dp_sink.vhd:363:34  */
  assign n13430_o = wr_burstlen_in[14:10];
  /* ../../HW/src/dp/dp_sink.vhd:364:30  */
  assign n13431_o = wr_bus_id_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:365:30  */
  assign n13432_o = wr_thread_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:366:36  */
  assign n13433_o = wr_data_type_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:367:38  */
  assign n13434_o = wr_data_model_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:368:28  */
  assign n13435_o = wr_mcast_in[17:12];
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13436_o = n13399_o ? n13402_o : n13420_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13437_o = n13399_o ? n13404_o : n13422_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13438_o = n13399_o ? n13405_o : n13423_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13439_o = n13399_o ? n13403_o : n13421_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13440_o = n13399_o ? n13406_o : n13424_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13441_o = n13399_o ? n13407_o : n13425_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13442_o = n13399_o ? n13408_o : n13426_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13443_o = n13399_o ? n13409_o : n13427_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13444_o = n13399_o ? n13410_o : n13428_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13445_o = n13399_o ? n13411_o : n13429_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13446_o = n13399_o ? n13400_o : n13418_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13447_o = n13399_o ? n13401_o : n13419_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13448_o = n13399_o ? n13412_o : n13430_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13449_o = n13399_o ? n13413_o : n13431_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13450_o = n13399_o ? n13414_o : n13432_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13451_o = n13399_o ? n13415_o : n13433_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13452_o = n13399_o ? n13416_o : n13434_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n13453_o = n13399_o ? n13417_o : n13435_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13454_o = n13380_o ? n13383_o : n13436_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13455_o = n13380_o ? n13385_o : n13437_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13456_o = n13380_o ? n13386_o : n13438_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13457_o = n13380_o ? n13384_o : n13439_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13458_o = n13380_o ? n13387_o : n13440_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13459_o = n13380_o ? n13388_o : n13441_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13460_o = n13380_o ? n13389_o : n13442_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13461_o = n13380_o ? n13390_o : n13443_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13462_o = n13380_o ? n13391_o : n13444_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13463_o = n13380_o ? n13392_o : n13445_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13464_o = n13380_o ? n13381_o : n13446_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13465_o = n13380_o ? n13382_o : n13447_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13466_o = n13380_o ? n13393_o : n13448_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13467_o = n13380_o ? n13394_o : n13449_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13468_o = n13380_o ? n13395_o : n13450_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13469_o = n13380_o ? n13396_o : n13451_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13470_o = n13380_o ? n13397_o : n13452_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n13471_o = n13380_o ? n13398_o : n13453_o;
  /* ../../HW/src/dp/dp_sink.vhd:464:17  */
  assign n13513_o = ~reset_in;
  /* ../../HW/src/dp/dp_sink.vhd:515:26  */
  assign n13516_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:515:53  */
  assign n13517_o = wr_datavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:515:34  */
  assign n13518_o = n13517_o & n13516_o;
  /* ../../HW/src/dp/dp_sink.vhd:515:70  */
  assign n13519_o = ~wr_vm;
  /* ../../HW/src/dp/dp_sink.vhd:515:61  */
  assign n13520_o = n13519_o & n13518_o;
  /* ../../HW/src/dp/dp_sink.vhd:516:41  */
  assign n13522_o = req_p0_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:515:13  */
  assign n13523_o = n13520_o ? n13522_o : req_p0_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:520:26  */
  assign n13524_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:520:53  */
  assign n13525_o = wr_datavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:520:34  */
  assign n13526_o = n13525_o & n13524_o;
  /* ../../HW/src/dp/dp_sink.vhd:520:70  */
  assign n13527_o = ~wr_vm;
  /* ../../HW/src/dp/dp_sink.vhd:520:61  */
  assign n13528_o = n13527_o & n13526_o;
  /* ../../HW/src/dp/dp_sink.vhd:521:41  */
  assign n13530_o = req_p0_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:520:13  */
  assign n13531_o = n13528_o ? n13530_o : req_p0_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:525:26  */
  assign n13532_o = wr_req_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:525:53  */
  assign n13533_o = wr_datavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:525:34  */
  assign n13534_o = n13533_o & n13532_o;
  /* ../../HW/src/dp/dp_sink.vhd:525:70  */
  assign n13535_o = ~wr_vm;
  /* ../../HW/src/dp/dp_sink.vhd:525:61  */
  assign n13536_o = n13535_o & n13534_o;
  /* ../../HW/src/dp/dp_sink.vhd:526:41  */
  assign n13538_o = req_p0_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:525:13  */
  assign n13539_o = n13536_o ? n13538_o : req_p0_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:533:26  */
  assign n13540_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:533:53  */
  assign n13541_o = wr_datavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:533:34  */
  assign n13542_o = n13541_o & n13540_o;
  /* ../../HW/src/dp/dp_sink.vhd:533:61  */
  assign n13543_o = wr_vm & n13542_o;
  /* ../../HW/src/dp/dp_sink.vhd:534:41  */
  assign n13545_o = req_p1_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:533:13  */
  assign n13546_o = n13543_o ? n13545_o : req_p1_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:538:26  */
  assign n13547_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:538:53  */
  assign n13548_o = wr_datavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:538:34  */
  assign n13549_o = n13548_o & n13547_o;
  /* ../../HW/src/dp/dp_sink.vhd:538:61  */
  assign n13550_o = wr_vm & n13549_o;
  /* ../../HW/src/dp/dp_sink.vhd:539:41  */
  assign n13552_o = req_p1_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:538:13  */
  assign n13553_o = n13550_o ? n13552_o : req_p1_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:543:26  */
  assign n13554_o = wr_req_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:543:53  */
  assign n13555_o = wr_datavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:543:34  */
  assign n13556_o = n13555_o & n13554_o;
  /* ../../HW/src/dp/dp_sink.vhd:543:61  */
  assign n13557_o = wr_vm & n13556_o;
  /* ../../HW/src/dp/dp_sink.vhd:544:41  */
  assign n13559_o = req_p1_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:543:13  */
  assign n13560_o = n13557_o ? n13559_o : req_p1_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:551:23  */
  assign n13561_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:551:57  */
  assign n13562_o = wr_readdatavalid_vm_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:551:60  */
  assign n13563_o = ~n13562_o;
  /* ../../HW/src/dp/dp_sink.vhd:551:31  */
  assign n13564_o = n13563_o & n13561_o;
  /* ../../HW/src/dp/dp_sink.vhd:552:41  */
  assign n13566_o = rsp_p0_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:551:13  */
  assign n13567_o = n13564_o ? n13566_o : rsp_p0_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:556:23  */
  assign n13568_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:556:57  */
  assign n13569_o = wr_readdatavalid_vm_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:556:60  */
  assign n13570_o = ~n13569_o;
  /* ../../HW/src/dp/dp_sink.vhd:556:31  */
  assign n13571_o = n13570_o & n13568_o;
  /* ../../HW/src/dp/dp_sink.vhd:557:41  */
  assign n13573_o = rsp_p0_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:556:13  */
  assign n13574_o = n13571_o ? n13573_o : rsp_p0_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:561:23  */
  assign n13575_o = wr_req2[2];
  /* ../../HW/src/dp/dp_sink.vhd:561:57  */
  assign n13576_o = wr_readdatavalid_vm_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:561:60  */
  assign n13577_o = ~n13576_o;
  /* ../../HW/src/dp/dp_sink.vhd:561:31  */
  assign n13578_o = n13577_o & n13575_o;
  /* ../../HW/src/dp/dp_sink.vhd:562:41  */
  assign n13580_o = rsp_p0_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:561:13  */
  assign n13581_o = n13578_o ? n13580_o : rsp_p0_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:569:23  */
  assign n13582_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:569:57  */
  assign n13583_o = wr_readdatavalid_vm_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:569:31  */
  assign n13584_o = n13583_o & n13582_o;
  /* ../../HW/src/dp/dp_sink.vhd:570:41  */
  assign n13586_o = rsp_p1_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:569:13  */
  assign n13587_o = n13584_o ? n13586_o : rsp_p1_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:574:23  */
  assign n13588_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:574:57  */
  assign n13589_o = wr_readdatavalid_vm_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:574:31  */
  assign n13590_o = n13589_o & n13588_o;
  /* ../../HW/src/dp/dp_sink.vhd:575:41  */
  assign n13592_o = rsp_p1_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:574:13  */
  assign n13593_o = n13590_o ? n13592_o : rsp_p1_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:579:23  */
  assign n13594_o = wr_req2[2];
  /* ../../HW/src/dp/dp_sink.vhd:579:57  */
  assign n13595_o = wr_readdatavalid_vm_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:579:31  */
  assign n13596_o = n13595_o & n13594_o;
  /* ../../HW/src/dp/dp_sink.vhd:580:41  */
  assign n13598_o = rsp_p1_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:579:13  */
  assign n13599_o = n13596_o ? n13598_o : rsp_p1_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:601:28  */
  assign n13600_o = n13523_o != n13567_o;
  /* ../../HW/src/dp/dp_sink.vhd:601:13  */
  assign n13603_o = n13600_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:607:28  */
  assign n13604_o = n13531_o != n13574_o;
  /* ../../HW/src/dp/dp_sink.vhd:607:13  */
  assign n13607_o = n13604_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:613:28  */
  assign n13608_o = n13539_o != n13581_o;
  /* ../../HW/src/dp/dp_sink.vhd:613:13  */
  assign n13611_o = n13608_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:621:28  */
  assign n13612_o = n13546_o != n13587_o;
  /* ../../HW/src/dp/dp_sink.vhd:621:13  */
  assign n13615_o = n13612_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:627:28  */
  assign n13616_o = n13553_o != n13593_o;
  /* ../../HW/src/dp/dp_sink.vhd:627:13  */
  assign n13619_o = n13616_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:633:28  */
  assign n13620_o = n13560_o != n13599_o;
  /* ../../HW/src/dp/dp_sink.vhd:633:13  */
  assign n13623_o = n13620_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:639:35  */
  assign n13624_o = ~bus_wait_request_in;
  /* ../../HW/src/dp/dp_sink.vhd:639:51  */
  assign n13625_o = ~valid_rr;
  /* ../../HW/src/dp/dp_sink.vhd:639:40  */
  assign n13626_o = n13624_o | n13625_o;
  /* ../../HW/src/dp/dp_sink.vhd:647:23  */
  assign n13627_o = q_r[0];
  /* ../../HW/src/dp/dp_sink.vhd:651:98  */
  assign n13628_o = q_r[64:1];
  /* ../../HW/src/dp/dp_sink.vhd:647:17  */
  assign n13629_o = n13627_o ? q2 : n13628_o;
  /* ../../HW/src/dp/dp_sink.vhd:656:49  */
  assign n13630_o = q_r[96:65];
  /* ../../HW/src/dp/dp_sink.vhd:659:34  */
  assign n13631_o = q_r[97];
  /* ../../HW/src/dp/dp_sink.vhd:661:39  */
  assign n13632_o = q_r[98];
  /* ../../HW/src/dp/dp_sink.vhd:663:32  */
  assign n13633_o = q_r[99];
  /* ../../HW/src/dp/dp_sink.vhd:666:51  */
  assign n13634_o = q_r[104:100];
  /* ../../HW/src/dp/dp_sink.vhd:667:27  */
  assign n13635_o = q_r[0];
  /* ../../HW/src/dp/dp_sink.vhd:668:52  */
  assign n13637_o = usedw2 + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:670:51  */
  assign n13639_o = usedw + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:667:21  */
  assign n13640_o = n13635_o ? n13637_o : n13639_o;
  assign n13642_o = {4'b0000, n13634_o};
  /* ../../HW/src/dp/dp_sink.vhd:674:31  */
  assign n13643_o = $unsigned(n13642_o) > $unsigned(n13640_o);
  /* ../../HW/src/dp/dp_sink.vhd:675:50  */
  assign n13644_o = n13640_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:674:21  */
  assign n13645_o = n13643_o ? n13644_o : n13634_o;
  /* ../../HW/src/dp/dp_sink.vhd:681:41  */
  assign n13646_o = q_r[106:105];
  /* ../../HW/src/dp/dp_sink.vhd:683:45  */
  assign n13647_o = q_r[107];
  /* ../../HW/src/dp/dp_sink.vhd:685:48  */
  assign n13648_o = q_r[109:108];
  /* ../../HW/src/dp/dp_sink.vhd:687:40  */
  assign n13649_o = q_r[111:110];
  /* ../../HW/src/dp/dp_sink.vhd:689:52  */
  assign n13650_o = q_r[117:112];
  /* ../../HW/src/dp/dp_sink.vhd:691:32  */
  assign n13651_o = q_r[120:118];
  /* ../../HW/src/dp/dp_sink.vhd:693:32  */
  assign n13652_o = q_r[121];
  /* ../../HW/src/dp/dp_sink.vhd:695:44  */
  assign n13653_o = q_r[123:122];
  /* ../../HW/src/dp/dp_sink.vhd:697:33  */
  assign n13654_o = q_r[125:124];
  /* ../../HW/src/dp/dp_sink.vhd:699:35  */
  assign n13655_o = q_r[127:126];
  /* ../../HW/src/dp/dp_sink.vhd:702:44  */
  assign n13656_o = q_r[131:128];
  /* ../../HW/src/dp/dp_sink.vhd:705:32  */
  assign n13657_o = {4'b0, n13645_o};  //  uext
  /* ../../HW/src/dp/dp_sink.vhd:706:38  */
  assign n13659_o = n13651_o == 3'b001;
  /* ../../HW/src/dp/dp_sink.vhd:707:35  */
  assign n13661_o = $unsigned(n13657_o) > $unsigned(9'b000010100);
  /* ../../HW/src/dp/dp_sink.vhd:707:20  */
  assign n13663_o = n13661_o ? 9'b000010011 : n13657_o;
  /* ../../HW/src/dp/dp_sink.vhd:710:50  */
  assign n13664_o = n13663_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:711:51  */
  assign n13666_o = n13663_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_sink.vhd:712:41  */
  assign n13668_o = n13651_o == 3'b011;
  /* ../../HW/src/dp/dp_sink.vhd:713:35  */
  assign n13670_o = $unsigned(n13657_o) > $unsigned(9'b000001010);
  /* ../../HW/src/dp/dp_sink.vhd:713:20  */
  assign n13672_o = n13670_o ? 9'b000001001 : n13657_o;
  /* ../../HW/src/dp/dp_sink.vhd:716:50  */
  assign n13673_o = n13672_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:717:51  */
  assign n13675_o = n13672_o << 32'b00000000000000000000000000000010;
  /* ../../HW/src/dp/dp_sink.vhd:718:41  */
  assign n13677_o = n13651_o == 3'b111;
  /* ../../HW/src/dp/dp_sink.vhd:719:35  */
  assign n13679_o = $unsigned(n13657_o) > $unsigned(9'b000000101);
  /* ../../HW/src/dp/dp_sink.vhd:719:20  */
  assign n13681_o = n13679_o ? 9'b000000100 : n13657_o;
  /* ../../HW/src/dp/dp_sink.vhd:722:50  */
  assign n13682_o = n13681_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:723:51  */
  assign n13684_o = n13681_o << 32'b00000000000000000000000000000011;
  /* ../../HW/src/dp/dp_sink.vhd:725:35  */
  assign n13686_o = $unsigned(n13657_o) > $unsigned(9'b000101000);
  /* ../../HW/src/dp/dp_sink.vhd:725:20  */
  assign n13688_o = n13686_o ? 9'b000100111 : n13657_o;
  /* ../../HW/src/dp/dp_sink.vhd:728:50  */
  assign n13689_o = n13688_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:718:17  */
  assign n13690_o = n13677_o ? n13684_o : n13688_o;
  /* ../../HW/src/dp/dp_sink.vhd:718:17  */
  assign n13691_o = n13677_o ? n13682_o : n13689_o;
  /* ../../HW/src/dp/dp_sink.vhd:712:17  */
  assign n13693_o = n13668_o ? n13675_o : n13690_o;
  /* ../../HW/src/dp/dp_sink.vhd:712:17  */
  assign n13694_o = n13668_o ? n13673_o : n13691_o;
  /* ../../HW/src/dp/dp_sink.vhd:706:17  */
  assign n13696_o = n13659_o ? n13666_o : n13693_o;
  /* ../../HW/src/dp/dp_sink.vhd:706:17  */
  assign n13697_o = n13659_o ? n13664_o : n13694_o;
  assign n13777_o = {n13611_o, n13607_o, n13603_o};
  assign n13779_o = {n13623_o, n13619_o, n13615_o};
  /* ../../HW/src/dp/dp_sink.vhd:759:12  */
  assign n14050_o = ~reset_in;
  /* ../../HW/src/dp/dp_sink.vhd:764:27  */
  assign n14052_o = ~usedw;
  /* ../../HW/src/dp/dp_sink.vhd:765:18  */
  assign n14054_o = $unsigned(n14052_o) <= $unsigned(9'b000101111);
  /* ../../HW/src/dp/dp_sink.vhd:765:7  */
  assign n14057_o = n14054_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:775:26  */
  assign n14072_o = ~empty;
  /* ../../HW/src/dp/dp_sink.vhd:775:44  */
  assign n14073_o = ~empty2;
  /* ../../HW/src/dp/dp_sink.vhd:775:54  */
  assign n14074_o = q[0];
  /* ../../HW/src/dp/dp_sink.vhd:775:57  */
  assign n14075_o = ~n14074_o;
  /* ../../HW/src/dp/dp_sink.vhd:775:50  */
  assign n14076_o = n14073_o | n14075_o;
  /* ../../HW/src/dp/dp_sink.vhd:775:32  */
  assign n14077_o = n14076_o & n14072_o;
  /* ../../HW/src/dp/dp_sink.vhd:775:15  */
  assign n14078_o = n14077_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:787:20  */
  assign n14082_o = q[0];
  /* ../../HW/src/dp/dp_sink.vhd:784:5  */
  assign n14084_o = emptyn ? emptyn : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:784:5  */
  assign n14086_o = emptyn ? n14082_o : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:784:5  */
  assign n14089_o = emptyn ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:780:5  */
  assign n14091_o = bus_wait_request_in ? 1'b0 : n14084_o;
  /* ../../HW/src/dp/dp_sink.vhd:780:5  */
  assign n14093_o = bus_wait_request_in ? 1'b0 : n14086_o;
  /* ../../HW/src/dp/dp_sink.vhd:780:5  */
  assign n14094_o = bus_wait_request_in ? valid_r : n14089_o;
  /* ../../HW/src/dp/dp_sink.vhd:797:20  */
  assign n14095_o = q[0];
  /* ../../HW/src/dp/dp_sink.vhd:794:5  */
  assign n14097_o = emptyn ? emptyn : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:794:5  */
  assign n14099_o = emptyn ? n14095_o : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:794:5  */
  assign n14102_o = emptyn ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:779:1  */
  assign n14103_o = valid_rr ? n14091_o : n14097_o;
  /* ../../HW/src/dp/dp_sink.vhd:779:1  */
  assign n14104_o = valid_rr ? n14093_o : n14099_o;
  /* ../../HW/src/dp/dp_sink.vhd:779:1  */
  assign n14105_o = valid_rr ? n14094_o : n14102_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14109_o = rdreq ? q : q_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14110_q <= 132'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n14110_q <= n14109_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14111_o = n13626_o ? valid : valid_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14112_q <= 1'b0;
    else
      n14112_q <= n14111_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14113_o = n13626_o ? valid_r : valid_rr;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14114_q <= 1'b0;
    else
      n14114_q <= n14113_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14115_o = n13626_o ? n13655_o : bus_data_flow_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14116_q <= 2'b00;
    else
      n14116_q <= n14115_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14117_o = n13626_o ? n13656_o : bus_end_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14118_q <= 4'b0000;
    else
      n14118_q <= n14117_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14119_o = n13626_o ? n13651_o : bus_vector_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14120_q <= 3'b000;
    else
      n14120_q <= n14119_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14121_o = n13626_o ? n13652_o : bus_stream_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14122_q <= 1'b0;
    else
      n14122_q <= n14121_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14123_o = n13626_o ? n13653_o : bus_stream_id_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14124_q <= 2'b00;
    else
      n14124_q <= n14123_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14125_o = n13626_o ? n13654_o : bus_scatter_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14126_q <= 2'b00;
    else
      n14126_q <= n14125_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14127_o = n13626_o ? n13630_o : bus_addr_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14128_q <= 32'b00000000000000000000000000000000;
    else
      n14128_q <= n14127_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14129_o = n13626_o ? n13631_o : bus_fork_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14130_q <= 1'b0;
    else
      n14130_q <= n14129_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14131_o = n13626_o ? n13632_o : bus_addr_mode_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14132_q <= 1'b0;
    else
      n14132_q <= n14131_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14133_o = n13626_o ? n13633_o : bus_vm_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14134_q <= 1'b0;
    else
      n14134_q <= n14133_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14135_o = n13626_o ? n13629_o : bus_writedata_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14136_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n14136_q <= n14135_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14137_o = n13626_o ? n13645_o : bus_burstlen_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14138_q <= 5'b00000;
    else
      n14138_q <= n14137_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14139_o = n13626_o ? n13696_o : bus_burstlen2_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14140_q <= 9'b000000000;
    else
      n14140_q <= n14139_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14141_o = n13626_o ? n13697_o : bus_burstlen3_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14142_q <= 5'b00000;
    else
      n14142_q <= n14141_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14143_o = n13626_o ? n13646_o : bus_id_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14144_q <= 2'b00;
    else
      n14144_q <= n14143_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14145_o = n13626_o ? n13647_o : bus_thread_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14146_q <= 1'b0;
    else
      n14146_q <= n14145_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14147_o = n13626_o ? n13648_o : bus_data_type_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14148_q <= 2'b00;
    else
      n14148_q <= n14147_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14149_o = n13626_o ? n13649_o : bus_data_model_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14150_q <= 2'b00;
    else
      n14150_q <= n14149_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n14151_o = n13626_o ? n13650_o : bus_mcast_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14152_q <= 6'b111111;
    else
      n14152_q <= n14151_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14153_q <= 9'b000000000;
    else
      n14153_q <= n13523_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14154_q <= 9'b000000000;
    else
      n14154_q <= n13531_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14155_q <= 9'b000000000;
    else
      n14155_q <= n13539_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14156_q <= 9'b000000000;
    else
      n14156_q <= n13567_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14157_q <= 9'b000000000;
    else
      n14157_q <= n13574_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14158_q <= 9'b000000000;
    else
      n14158_q <= n13581_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14159_q <= 9'b000000000;
    else
      n14159_q <= n13546_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14160_q <= 9'b000000000;
    else
      n14160_q <= n13553_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14161_q <= 9'b000000000;
    else
      n14161_q <= n13560_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14162_q <= 9'b000000000;
    else
      n14162_q <= n13587_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14163_q <= 9'b000000000;
    else
      n14163_q <= n13593_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14164_q <= 9'b000000000;
    else
      n14164_q <= n13599_o;
  /* ../../HW/src/dp/dp_sink.vhd:464:5  */
  assign n14165_o = {wr_end, wr_data_flow, wr_scatter, wr_stream_id, wr_stream, wr_vector, wr_mcast, wr_data_model, wr_data_type, wr_thread, wr_bus_id, wr_burstlen, wr_vm, wr_addr_mode, wr_fork, wr_addr, wr_data, wr_datavalid};
  /* ../../HW/src/dp/dp_sink.vhd:464:5  */
  assign n14166_o = {n13359_o, n13351_o, n13343_o};
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14167_q <= 3'b000;
    else
      n14167_q <= n13777_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n13513_o)
    if (n13513_o)
      n14168_q <= 3'b000;
    else
      n14168_q <= n13779_o;
  /* ../../HW/src/dp/dp_sink.vhd:763:4  */
  always @(posedge clock_in or posedge n14050_o)
    if (n14050_o)
      n14169_q <= 1'b0;
    else
      n14169_q <= n14057_o;
  /* ../../HW/src/dp/dp_sink.vhd:763:4  */
  always @(posedge clock_in or posedge n14050_o)
    if (n14050_o)
      n14170_q <= 5'b00000;
    else
      n14170_q <= 5'b11111;
endmodule

module dp_sink_3_32_1_9_6a0e3f59309a30c5143aeb870000c064ad45653d
  (input  clock_in,
   input  reset_in,
   input  bus_wait_request_in,
   input  [2:0] wr_req_in,
   input  [2:0] wr_req_pending_p0_in,
   input  [2:0] wr_req_pending_p1_in,
   input  [5:0] wr_data_flow_in,
   input  [8:0] wr_vector_in,
   input  [2:0] wr_stream_in,
   input  [5:0] wr_stream_id_in,
   input  [5:0] wr_scatter_in,
   input  [11:0] wr_end_in,
   input  [95:0] wr_addr_in,
   input  [2:0] wr_fork_in,
   input  [2:0] wr_addr_mode_in,
   input  [2:0] wr_src_vm_in,
   input  [2:0] wr_datavalid_in,
   input  [191:0] wr_data_in,
   input  [2:0] wr_readdatavalid_in,
   input  [2:0] wr_readdatavalid_vm_in,
   input  [191:0] wr_readdata_in,
   input  [14:0] wr_burstlen_in,
   input  [5:0] wr_bus_id_in,
   input  [2:0] wr_thread_in,
   input  [5:0] wr_data_type_in,
   input  [5:0] wr_data_model_in,
   input  [17:0] wr_mcast_in,
   output [31:0] bus_addr_out,
   output bus_fork_out,
   output bus_addr_mode_out,
   output bus_vm_out,
   output [1:0] bus_data_flow_out,
   output [2:0] bus_vector_out,
   output bus_stream_out,
   output [1:0] bus_stream_id_out,
   output [1:0] bus_scatter_out,
   output [3:0] bus_end_out,
   output [5:0] bus_mcast_out,
   output bus_cs_out,
   output bus_write_out,
   output [63:0] bus_writedata_out,
   output [4:0] bus_burstlen_out,
   output [8:0] bus_burstlen2_out,
   output [4:0] bus_burstlen3_out,
   output [1:0] bus_id_out,
   output [1:0] bus_data_type_out,
   output [1:0] bus_data_model_out,
   output bus_thread_out,
   output [4:0] wr_maxburstlen_out,
   output wr_full_out,
   output [2:0] read_pending_p0_out,
   output [2:0] read_pending_p1_out);
  wire rdreq;
  wire rdreq2;
  wire empty;
  wire emptyn;
  wire empty2;
  wire [63:0] q2;
  wire [131:0] q;
  wire [131:0] q_r;
  wire valid;
  wire valid_r;
  wire valid_rr;
  wire [1:0] bus_data_flow_r;
  wire [3:0] bus_end_r;
  wire [2:0] bus_vector_r;
  wire bus_stream_r;
  wire [1:0] bus_stream_id_r;
  wire [1:0] bus_scatter_r;
  wire [31:0] bus_addr_r;
  wire bus_fork_r;
  wire bus_addr_mode_r;
  wire bus_vm_r;
  wire [63:0] bus_writedata_r;
  wire [4:0] bus_burstlen_r;
  wire [8:0] bus_burstlen2_r;
  wire [4:0] bus_burstlen3_r;
  wire [1:0] bus_id_r;
  wire bus_thread_r;
  wire [1:0] bus_data_type_r;
  wire [1:0] bus_data_model_r;
  reg [5:0] bus_mcast_r;
  wire [8:0] req_p0_0_r;
  wire [8:0] req_p0_1_r;
  wire [8:0] req_p0_2_r;
  wire [8:0] rsp_p0_0_r;
  wire [8:0] rsp_p0_1_r;
  wire [8:0] rsp_p0_2_r;
  wire [8:0] req_p1_0_r;
  wire [8:0] req_p1_1_r;
  wire [8:0] req_p1_2_r;
  wire [8:0] rsp_p1_0_r;
  wire [8:0] rsp_p1_1_r;
  wire [8:0] rsp_p1_2_r;
  wire [8:0] usedw;
  wire [131:0] fifo_data;
  wire [31:0] wr_addr;
  wire wr_fork;
  wire wr_addr_mode;
  wire wr_vm;
  wire [1:0] wr_data_flow;
  wire [2:0] wr_vector;
  wire wr_stream;
  wire [1:0] wr_stream_id;
  wire [1:0] wr_scatter;
  wire [3:0] wr_end;
  wire wr_datavalid;
  wire [63:0] wr_data;
  wire [63:0] wr_data2;
  wire [4:0] wr_burstlen;
  wire [1:0] wr_bus_id;
  wire wr_thread;
  wire [1:0] wr_data_type;
  wire [1:0] wr_data_model;
  wire [5:0] wr_mcast;
  wire wr_req;
  wire [2:0] wr_req2;
  wire wr_req2_all;
  wire [2:0] read_pending_p0_r;
  wire [2:0] read_pending_p1_r;
  wire wr_full_r;
  wire [4:0] wr_maxburstlen_r;
  wire [131:0] dp_sink_fifo_i_n12425;
  wire [8:0] dp_sink_fifo_i_n12427;
  wire dp_sink_fifo_i_n12428;
  wire [131:0] dp_sink_fifo_i_q_out;
  wire [8:0] dp_sink_fifo_i_ravail_out;
  wire [8:0] dp_sink_fifo_i_wused_out;
  wire dp_sink_fifo_i_empty_out;
  wire dp_sink_fifo_i_full_out;
  wire dp_sink_fifo_i_almost_full_out;
  wire [63:0] dp_sink_fifo_i2_n12441;
  wire dp_sink_fifo_i2_n12444;
  wire [63:0] dp_sink_fifo_i2_q_out;
  wire [8:0] dp_sink_fifo_i2_ravail_out;
  wire [8:0] dp_sink_fifo_i2_wused_out;
  wire dp_sink_fifo_i2_empty_out;
  wire dp_sink_fifo_i2_full_out;
  wire dp_sink_fifo_i2_almost_full_out;
  wire n12457_o;
  wire n12458_o;
  wire n12459_o;
  wire n12460_o;
  wire n12461_o;
  wire n12463_o;
  wire n12464_o;
  wire n12465_o;
  wire n12466_o;
  wire n12467_o;
  wire n12468_o;
  wire n12471_o;
  wire n12472_o;
  wire n12473_o;
  wire n12474_o;
  wire n12475_o;
  wire n12476_o;
  wire n12479_o;
  wire n12480_o;
  wire n12481_o;
  wire n12482_o;
  wire n12483_o;
  wire n12484_o;
  wire n12486_o;
  wire n12487_o;
  wire n12488_o;
  wire n12489_o;
  wire n12490_o;
  wire [2:0] n12491_o;
  wire [2:0] n12492_o;
  wire n12495_o;
  wire [63:0] n12496_o;
  wire n12497_o;
  wire [63:0] n12498_o;
  wire [63:0] n12499_o;
  wire [63:0] n12500_o;
  wire [63:0] n12501_o;
  wire n12505_o;
  wire n12506_o;
  wire [63:0] n12507_o;
  wire [31:0] n12508_o;
  wire n12509_o;
  wire n12510_o;
  wire n12511_o;
  wire [1:0] n12512_o;
  wire [2:0] n12513_o;
  wire n12514_o;
  wire [1:0] n12515_o;
  wire [1:0] n12516_o;
  wire [3:0] n12517_o;
  wire [4:0] n12518_o;
  wire [1:0] n12519_o;
  wire n12520_o;
  wire [1:0] n12521_o;
  wire [1:0] n12522_o;
  wire [5:0] n12523_o;
  wire n12524_o;
  wire n12525_o;
  wire [63:0] n12526_o;
  wire [31:0] n12527_o;
  wire n12528_o;
  wire n12529_o;
  wire n12530_o;
  wire [1:0] n12531_o;
  wire [2:0] n12532_o;
  wire n12533_o;
  wire [1:0] n12534_o;
  wire [1:0] n12535_o;
  wire [3:0] n12536_o;
  wire [4:0] n12537_o;
  wire [1:0] n12538_o;
  wire n12539_o;
  wire [1:0] n12540_o;
  wire [1:0] n12541_o;
  wire [5:0] n12542_o;
  wire n12543_o;
  wire [63:0] n12544_o;
  wire [31:0] n12545_o;
  wire n12546_o;
  wire n12547_o;
  wire n12548_o;
  wire [1:0] n12549_o;
  wire [2:0] n12550_o;
  wire n12551_o;
  wire [1:0] n12552_o;
  wire [1:0] n12553_o;
  wire [3:0] n12554_o;
  wire [4:0] n12555_o;
  wire [1:0] n12556_o;
  wire n12557_o;
  wire [1:0] n12558_o;
  wire [1:0] n12559_o;
  wire [5:0] n12560_o;
  wire [31:0] n12561_o;
  wire n12562_o;
  wire n12563_o;
  wire n12564_o;
  wire [1:0] n12565_o;
  wire [2:0] n12566_o;
  wire n12567_o;
  wire [1:0] n12568_o;
  wire [1:0] n12569_o;
  wire [3:0] n12570_o;
  wire n12571_o;
  wire [63:0] n12572_o;
  wire [4:0] n12573_o;
  wire [1:0] n12574_o;
  wire n12575_o;
  wire [1:0] n12576_o;
  wire [1:0] n12577_o;
  wire [5:0] n12578_o;
  wire [31:0] n12579_o;
  wire n12580_o;
  wire n12581_o;
  wire n12582_o;
  wire [1:0] n12583_o;
  wire [2:0] n12584_o;
  wire n12585_o;
  wire [1:0] n12586_o;
  wire [1:0] n12587_o;
  wire [3:0] n12588_o;
  wire n12589_o;
  wire [63:0] n12590_o;
  wire [4:0] n12591_o;
  wire [1:0] n12592_o;
  wire n12593_o;
  wire [1:0] n12594_o;
  wire [1:0] n12595_o;
  wire [5:0] n12596_o;
  wire n12638_o;
  wire n12641_o;
  wire n12642_o;
  wire n12643_o;
  wire n12644_o;
  wire n12645_o;
  wire [8:0] n12647_o;
  wire [8:0] n12648_o;
  wire n12649_o;
  wire n12650_o;
  wire n12651_o;
  wire n12652_o;
  wire n12653_o;
  wire [8:0] n12655_o;
  wire [8:0] n12656_o;
  wire n12657_o;
  wire n12658_o;
  wire n12659_o;
  wire n12660_o;
  wire n12661_o;
  wire [8:0] n12663_o;
  wire [8:0] n12664_o;
  wire n12665_o;
  wire n12666_o;
  wire n12667_o;
  wire n12668_o;
  wire [8:0] n12670_o;
  wire [8:0] n12671_o;
  wire n12672_o;
  wire n12673_o;
  wire n12674_o;
  wire n12675_o;
  wire [8:0] n12677_o;
  wire [8:0] n12678_o;
  wire n12679_o;
  wire n12680_o;
  wire n12681_o;
  wire n12682_o;
  wire [8:0] n12684_o;
  wire [8:0] n12685_o;
  wire n12686_o;
  wire n12687_o;
  wire n12688_o;
  wire n12689_o;
  wire [8:0] n12691_o;
  wire [8:0] n12692_o;
  wire n12693_o;
  wire n12694_o;
  wire n12695_o;
  wire n12696_o;
  wire [8:0] n12698_o;
  wire [8:0] n12699_o;
  wire n12700_o;
  wire n12701_o;
  wire n12702_o;
  wire n12703_o;
  wire [8:0] n12705_o;
  wire [8:0] n12706_o;
  wire n12707_o;
  wire n12708_o;
  wire n12709_o;
  wire [8:0] n12711_o;
  wire [8:0] n12712_o;
  wire n12713_o;
  wire n12714_o;
  wire n12715_o;
  wire [8:0] n12717_o;
  wire [8:0] n12718_o;
  wire n12719_o;
  wire n12720_o;
  wire n12721_o;
  wire [8:0] n12723_o;
  wire [8:0] n12724_o;
  wire n12725_o;
  wire n12728_o;
  wire n12729_o;
  wire n12732_o;
  wire n12733_o;
  wire n12736_o;
  wire n12737_o;
  wire n12740_o;
  wire n12741_o;
  wire n12744_o;
  wire n12745_o;
  wire n12748_o;
  wire n12749_o;
  wire n12750_o;
  wire n12751_o;
  wire n12752_o;
  wire [63:0] n12753_o;
  wire [63:0] n12754_o;
  wire [31:0] n12755_o;
  wire n12756_o;
  wire n12757_o;
  wire n12758_o;
  wire [1:0] n12759_o;
  wire n12760_o;
  wire [1:0] n12761_o;
  wire [1:0] n12762_o;
  wire [5:0] n12763_o;
  wire [2:0] n12764_o;
  wire n12765_o;
  wire [1:0] n12766_o;
  wire [1:0] n12767_o;
  wire [1:0] n12768_o;
  wire [3:0] n12769_o;
  wire n12773_o;
  wire n12775_o;
  wire [8:0] n12777_o;
  wire [4:0] n12778_o;
  wire [8:0] n12780_o;
  wire n12782_o;
  wire n12784_o;
  wire [8:0] n12786_o;
  wire [4:0] n12787_o;
  wire [8:0] n12789_o;
  wire n12791_o;
  wire n12793_o;
  wire [8:0] n12795_o;
  wire [4:0] n12796_o;
  wire [8:0] n12798_o;
  wire n12800_o;
  wire [8:0] n12802_o;
  wire [4:0] n12803_o;
  wire [8:0] n12804_o;
  wire [4:0] n12805_o;
  wire [8:0] n12807_o;
  wire [4:0] n12808_o;
  wire [8:0] n12810_o;
  wire [4:0] n12811_o;
  wire [2:0] n12890_o;
  wire [2:0] n12892_o;
  wire n13151_o;
  wire [8:0] n13153_o;
  wire n13155_o;
  wire n13158_o;
  wire n13173_o;
  wire n13174_o;
  wire n13175_o;
  wire n13176_o;
  wire n13177_o;
  wire n13178_o;
  wire n13179_o;
  wire n13183_o;
  wire n13185_o;
  wire n13187_o;
  wire n13190_o;
  wire n13192_o;
  wire n13194_o;
  wire n13195_o;
  wire n13196_o;
  wire n13198_o;
  wire n13200_o;
  wire n13203_o;
  wire n13204_o;
  wire n13205_o;
  wire n13206_o;
  wire [131:0] n13210_o;
  reg [131:0] n13211_q;
  wire n13212_o;
  reg n13213_q;
  wire n13214_o;
  reg n13215_q;
  wire [1:0] n13216_o;
  reg [1:0] n13217_q;
  wire [3:0] n13218_o;
  reg [3:0] n13219_q;
  wire [2:0] n13220_o;
  reg [2:0] n13221_q;
  wire n13222_o;
  reg n13223_q;
  wire [1:0] n13224_o;
  reg [1:0] n13225_q;
  wire [1:0] n13226_o;
  reg [1:0] n13227_q;
  wire [31:0] n13228_o;
  reg [31:0] n13229_q;
  wire n13230_o;
  reg n13231_q;
  wire n13232_o;
  reg n13233_q;
  wire n13234_o;
  reg n13235_q;
  wire [63:0] n13236_o;
  reg [63:0] n13237_q;
  wire [4:0] n13238_o;
  reg [4:0] n13239_q;
  wire [8:0] n13240_o;
  reg [8:0] n13241_q;
  wire [4:0] n13242_o;
  reg [4:0] n13243_q;
  wire [1:0] n13244_o;
  reg [1:0] n13245_q;
  wire n13246_o;
  reg n13247_q;
  wire [1:0] n13248_o;
  reg [1:0] n13249_q;
  wire [1:0] n13250_o;
  reg [1:0] n13251_q;
  wire [5:0] n13252_o;
  reg [5:0] n13253_q;
  reg [8:0] n13254_q;
  reg [8:0] n13255_q;
  reg [8:0] n13256_q;
  reg [8:0] n13257_q;
  reg [8:0] n13258_q;
  reg [8:0] n13259_q;
  reg [8:0] n13260_q;
  reg [8:0] n13261_q;
  reg [8:0] n13262_q;
  reg [8:0] n13263_q;
  reg [8:0] n13264_q;
  reg [8:0] n13265_q;
  wire [131:0] n13266_o;
  wire [2:0] n13267_o;
  reg [2:0] n13268_q;
  reg [2:0] n13269_q;
  reg n13270_q;
  reg [4:0] n13271_q;
  assign bus_addr_out = bus_addr_r;
  assign bus_fork_out = bus_fork_r;
  assign bus_addr_mode_out = bus_addr_mode_r;
  assign bus_vm_out = bus_vm_r;
  assign bus_data_flow_out = bus_data_flow_r;
  assign bus_vector_out = bus_vector_r;
  assign bus_stream_out = bus_stream_r;
  assign bus_stream_id_out = bus_stream_id_r;
  assign bus_scatter_out = bus_scatter_r;
  assign bus_end_out = bus_end_r;
  assign bus_mcast_out = bus_mcast_r;
  assign bus_cs_out = valid_rr;
  assign bus_write_out = valid_rr;
  assign bus_writedata_out = bus_writedata_r;
  assign bus_burstlen_out = bus_burstlen_r;
  assign bus_burstlen2_out = bus_burstlen2_r;
  assign bus_burstlen3_out = bus_burstlen3_r;
  assign bus_id_out = bus_id_r;
  assign bus_data_type_out = bus_data_type_r;
  assign bus_data_model_out = bus_data_model_r;
  assign bus_thread_out = bus_thread_r;
  assign wr_maxburstlen_out = wr_maxburstlen_r;
  assign wr_full_out = wr_full_r;
  assign read_pending_p0_out = n12491_o;
  assign read_pending_p1_out = n12492_o;
  /* ../../HW/src/dp/dp_sink.vhd:104:8  */
  assign rdreq = n13204_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:105:8  */
  assign rdreq2 = n13205_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:107:8  */
  assign empty = dp_sink_fifo_i_n12428; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:108:8  */
  assign emptyn = n13179_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:109:8  */
  assign empty2 = dp_sink_fifo_i2_n12444; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:110:8  */
  assign q2 = dp_sink_fifo_i2_n12441; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:113:8  */
  assign q = dp_sink_fifo_i_n12425; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:114:8  */
  assign q_r = n13211_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:115:8  */
  assign valid = n13206_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:116:8  */
  assign valid_r = n13213_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:117:8  */
  assign valid_rr = n13215_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:118:8  */
  assign bus_data_flow_r = n13217_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:119:8  */
  assign bus_end_r = n13219_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:120:8  */
  assign bus_vector_r = n13221_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:121:8  */
  assign bus_stream_r = n13223_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:122:8  */
  assign bus_stream_id_r = n13225_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:123:8  */
  assign bus_scatter_r = n13227_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:124:8  */
  assign bus_addr_r = n13229_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:125:8  */
  assign bus_fork_r = n13231_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:126:8  */
  assign bus_addr_mode_r = n13233_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:127:8  */
  assign bus_vm_r = n13235_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:128:8  */
  assign bus_writedata_r = n13237_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:129:8  */
  assign bus_burstlen_r = n13239_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:130:8  */
  assign bus_burstlen2_r = n13241_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:131:8  */
  assign bus_burstlen3_r = n13243_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:132:8  */
  assign bus_id_r = n13245_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:133:8  */
  assign bus_thread_r = n13247_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:134:8  */
  assign bus_data_type_r = n13249_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:135:8  */
  assign bus_data_model_r = n13251_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:136:8  */
  always @*
    bus_mcast_r = n13253_q; // (isignal)
  initial
    bus_mcast_r = 6'b111111;
  /* ../../HW/src/dp/dp_sink.vhd:137:8  */
  assign req_p0_0_r = n13254_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:138:8  */
  assign req_p0_1_r = n13255_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:139:8  */
  assign req_p0_2_r = n13256_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:140:8  */
  assign rsp_p0_0_r = n13257_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:141:8  */
  assign rsp_p0_1_r = n13258_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:142:8  */
  assign rsp_p0_2_r = n13259_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:144:8  */
  assign req_p1_0_r = n13260_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:145:8  */
  assign req_p1_1_r = n13261_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:146:8  */
  assign req_p1_2_r = n13262_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:147:8  */
  assign rsp_p1_0_r = n13263_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:148:8  */
  assign rsp_p1_1_r = n13264_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:149:8  */
  assign rsp_p1_2_r = n13265_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:155:8  */
  assign usedw = dp_sink_fifo_i_n12427; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:157:8  */
  assign fifo_data = n13266_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:159:8  */
  assign wr_addr = n12579_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:160:8  */
  assign wr_fork = n12580_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:161:8  */
  assign wr_addr_mode = n12581_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:162:8  */
  assign wr_vm = n12582_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:163:8  */
  assign wr_data_flow = n12583_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:164:8  */
  assign wr_vector = n12584_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:165:8  */
  assign wr_stream = n12585_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:166:8  */
  assign wr_stream_id = n12586_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:167:8  */
  assign wr_scatter = n12587_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:168:8  */
  assign wr_end = n12588_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:169:8  */
  assign wr_datavalid = n12589_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:170:8  */
  assign wr_data = n12590_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:171:8  */
  assign wr_data2 = n12501_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:172:8  */
  assign wr_burstlen = n12591_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:173:8  */
  assign wr_bus_id = n12592_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:174:8  */
  assign wr_thread = n12593_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:175:8  */
  assign wr_data_type = n12594_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:176:8  */
  assign wr_data_model = n12595_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:177:8  */
  assign wr_mcast = n12596_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:178:8  */
  assign wr_req = n12461_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:179:8  */
  assign wr_req2 = n13267_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:180:8  */
  assign wr_req2_all = n12490_o; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:185:8  */
  assign read_pending_p0_r = n13268_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:186:8  */
  assign read_pending_p1_r = n13269_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:188:8  */
  assign wr_full_r = n13270_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:189:8  */
  assign wr_maxburstlen_r = n13271_q; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:222:16  */
  assign dp_sink_fifo_i_n12425 = dp_sink_fifo_i_q_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:224:20  */
  assign dp_sink_fifo_i_n12427 = dp_sink_fifo_i_wused_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:225:20  */
  assign dp_sink_fifo_i_n12428 = dp_sink_fifo_i_empty_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:208:1  */
  scfifo_132_9_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 dp_sink_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(fifo_data),
    .write_in(wr_req),
    .read_in(rdreq),
    .q_out(dp_sink_fifo_i_q_out),
    .ravail_out(),
    .wused_out(dp_sink_fifo_i_wused_out),
    .empty_out(dp_sink_fifo_i_empty_out),
    .full_out(),
    .almost_full_out());
  /* ../../HW/src/dp/dp_sink.vhd:244:16  */
  assign dp_sink_fifo_i2_n12441 = dp_sink_fifo_i2_q_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:247:20  */
  assign dp_sink_fifo_i2_n12444 = dp_sink_fifo_i2_empty_out; // (signal)
  /* ../../HW/src/dp/dp_sink.vhd:230:1  */
  scfifo_64_9_1_5ba93c9db0cff93f52b521d7420e43f6eda2784f dp_sink_fifo_i2 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(wr_data2),
    .write_in(wr_req2_all),
    .read_in(rdreq2),
    .q_out(dp_sink_fifo_i2_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(dp_sink_fifo_i2_empty_out),
    .full_out(),
    .almost_full_out());
  /* ../../HW/src/dp/dp_sink.vhd:282:20  */
  assign n12457_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:282:36  */
  assign n12458_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:282:24  */
  assign n12459_o = n12457_o | n12458_o;
  /* ../../HW/src/dp/dp_sink.vhd:282:52  */
  assign n12460_o = wr_req_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:282:40  */
  assign n12461_o = n12459_o | n12460_o;
  /* ../../HW/src/dp/dp_sink.vhd:284:44  */
  assign n12463_o = wr_readdatavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:284:68  */
  assign n12464_o = req_p0_0_r != rsp_p0_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:284:96  */
  assign n12465_o = req_p1_0_r != rsp_p1_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:284:82  */
  assign n12466_o = n12464_o | n12465_o;
  /* ../../HW/src/dp/dp_sink.vhd:284:52  */
  assign n12467_o = n12466_o & n12463_o;
  /* ../../HW/src/dp/dp_sink.vhd:284:19  */
  assign n12468_o = n12467_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:286:44  */
  assign n12471_o = wr_readdatavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:286:68  */
  assign n12472_o = req_p0_1_r != rsp_p0_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:286:96  */
  assign n12473_o = req_p1_1_r != rsp_p1_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:286:82  */
  assign n12474_o = n12472_o | n12473_o;
  /* ../../HW/src/dp/dp_sink.vhd:286:52  */
  assign n12475_o = n12474_o & n12471_o;
  /* ../../HW/src/dp/dp_sink.vhd:286:19  */
  assign n12476_o = n12475_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:288:44  */
  assign n12479_o = wr_readdatavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:288:68  */
  assign n12480_o = req_p0_2_r != rsp_p0_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:288:96  */
  assign n12481_o = req_p1_2_r != rsp_p1_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:288:82  */
  assign n12482_o = n12480_o | n12481_o;
  /* ../../HW/src/dp/dp_sink.vhd:288:52  */
  assign n12483_o = n12482_o & n12479_o;
  /* ../../HW/src/dp/dp_sink.vhd:288:19  */
  assign n12484_o = n12483_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:290:23  */
  assign n12486_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:290:37  */
  assign n12487_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:290:27  */
  assign n12488_o = n12486_o | n12487_o;
  /* ../../HW/src/dp/dp_sink.vhd:290:51  */
  assign n12489_o = wr_req2[2];
  /* ../../HW/src/dp/dp_sink.vhd:290:41  */
  assign n12490_o = n12488_o | n12489_o;
  /* ../../HW/src/dp/dp_sink.vhd:292:42  */
  assign n12491_o = read_pending_p0_r | wr_req_pending_p0_in;
  /* ../../HW/src/dp/dp_sink.vhd:294:42  */
  assign n12492_o = read_pending_p1_r | wr_req_pending_p1_in;
  /* ../../HW/src/dp/dp_sink.vhd:299:14  */
  assign n12495_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:300:88  */
  assign n12496_o = wr_readdata_in[63:0];
  /* ../../HW/src/dp/dp_sink.vhd:301:17  */
  assign n12497_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:302:88  */
  assign n12498_o = wr_readdata_in[127:64];
  /* ../../HW/src/dp/dp_sink.vhd:304:88  */
  assign n12499_o = wr_readdata_in[191:128];
  /* ../../HW/src/dp/dp_sink.vhd:301:4  */
  assign n12500_o = n12497_o ? n12498_o : n12499_o;
  /* ../../HW/src/dp/dp_sink.vhd:299:4  */
  assign n12501_o = n12495_o ? n12496_o : n12500_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:13  */
  assign n12505_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:313:36  */
  assign n12506_o = wr_datavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:314:26  */
  assign n12507_o = wr_data_in[63:0];
  /* ../../HW/src/dp/dp_sink.vhd:315:26  */
  assign n12508_o = wr_addr_in[31:0];
  /* ../../HW/src/dp/dp_sink.vhd:316:26  */
  assign n12509_o = wr_src_vm_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:317:29  */
  assign n12510_o = wr_fork_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:318:36  */
  assign n12511_o = wr_addr_mode_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:319:36  */
  assign n12512_o = wr_data_flow_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:320:30  */
  assign n12513_o = wr_vector_in[2:0];
  /* ../../HW/src/dp/dp_sink.vhd:321:30  */
  assign n12514_o = wr_stream_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:322:36  */
  assign n12515_o = wr_stream_id_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:323:32  */
  assign n12516_o = wr_scatter_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:324:24  */
  assign n12517_o = wr_end_in[3:0];
  /* ../../HW/src/dp/dp_sink.vhd:325:34  */
  assign n12518_o = wr_burstlen_in[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:326:30  */
  assign n12519_o = wr_bus_id_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:327:30  */
  assign n12520_o = wr_thread_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:328:36  */
  assign n12521_o = wr_data_type_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:329:38  */
  assign n12522_o = wr_data_model_in[1:0];
  /* ../../HW/src/dp/dp_sink.vhd:330:28  */
  assign n12523_o = wr_mcast_in[5:0];
  /* ../../HW/src/dp/dp_sink.vhd:331:16  */
  assign n12524_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:332:36  */
  assign n12525_o = wr_datavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:333:26  */
  assign n12526_o = wr_data_in[127:64];
  /* ../../HW/src/dp/dp_sink.vhd:334:26  */
  assign n12527_o = wr_addr_in[63:32];
  /* ../../HW/src/dp/dp_sink.vhd:335:26  */
  assign n12528_o = wr_src_vm_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:336:29  */
  assign n12529_o = wr_fork_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:337:36  */
  assign n12530_o = wr_addr_mode_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:338:36  */
  assign n12531_o = wr_data_flow_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:339:30  */
  assign n12532_o = wr_vector_in[5:3];
  /* ../../HW/src/dp/dp_sink.vhd:340:30  */
  assign n12533_o = wr_stream_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:341:36  */
  assign n12534_o = wr_stream_id_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:342:32  */
  assign n12535_o = wr_scatter_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:343:24  */
  assign n12536_o = wr_end_in[7:4];
  /* ../../HW/src/dp/dp_sink.vhd:344:34  */
  assign n12537_o = wr_burstlen_in[9:5];
  /* ../../HW/src/dp/dp_sink.vhd:345:30  */
  assign n12538_o = wr_bus_id_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:346:30  */
  assign n12539_o = wr_thread_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:347:36  */
  assign n12540_o = wr_data_type_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:348:38  */
  assign n12541_o = wr_data_model_in[3:2];
  /* ../../HW/src/dp/dp_sink.vhd:349:28  */
  assign n12542_o = wr_mcast_in[11:6];
  /* ../../HW/src/dp/dp_sink.vhd:351:36  */
  assign n12543_o = wr_datavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:352:26  */
  assign n12544_o = wr_data_in[191:128];
  /* ../../HW/src/dp/dp_sink.vhd:353:26  */
  assign n12545_o = wr_addr_in[95:64];
  /* ../../HW/src/dp/dp_sink.vhd:354:26  */
  assign n12546_o = wr_src_vm_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:355:29  */
  assign n12547_o = wr_fork_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:356:36  */
  assign n12548_o = wr_addr_mode_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:357:36  */
  assign n12549_o = wr_data_flow_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:358:30  */
  assign n12550_o = wr_vector_in[8:6];
  /* ../../HW/src/dp/dp_sink.vhd:359:30  */
  assign n12551_o = wr_stream_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:360:36  */
  assign n12552_o = wr_stream_id_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:361:32  */
  assign n12553_o = wr_scatter_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:362:24  */
  assign n12554_o = wr_end_in[11:8];
  /* ../../HW/src/dp/dp_sink.vhd:363:34  */
  assign n12555_o = wr_burstlen_in[14:10];
  /* ../../HW/src/dp/dp_sink.vhd:364:30  */
  assign n12556_o = wr_bus_id_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:365:30  */
  assign n12557_o = wr_thread_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:366:36  */
  assign n12558_o = wr_data_type_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:367:38  */
  assign n12559_o = wr_data_model_in[5:4];
  /* ../../HW/src/dp/dp_sink.vhd:368:28  */
  assign n12560_o = wr_mcast_in[17:12];
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12561_o = n12524_o ? n12527_o : n12545_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12562_o = n12524_o ? n12529_o : n12547_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12563_o = n12524_o ? n12530_o : n12548_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12564_o = n12524_o ? n12528_o : n12546_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12565_o = n12524_o ? n12531_o : n12549_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12566_o = n12524_o ? n12532_o : n12550_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12567_o = n12524_o ? n12533_o : n12551_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12568_o = n12524_o ? n12534_o : n12552_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12569_o = n12524_o ? n12535_o : n12553_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12570_o = n12524_o ? n12536_o : n12554_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12571_o = n12524_o ? n12525_o : n12543_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12572_o = n12524_o ? n12526_o : n12544_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12573_o = n12524_o ? n12537_o : n12555_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12574_o = n12524_o ? n12538_o : n12556_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12575_o = n12524_o ? n12539_o : n12557_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12576_o = n12524_o ? n12540_o : n12558_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12577_o = n12524_o ? n12541_o : n12559_o;
  /* ../../HW/src/dp/dp_sink.vhd:331:1  */
  assign n12578_o = n12524_o ? n12542_o : n12560_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12579_o = n12505_o ? n12508_o : n12561_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12580_o = n12505_o ? n12510_o : n12562_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12581_o = n12505_o ? n12511_o : n12563_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12582_o = n12505_o ? n12509_o : n12564_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12583_o = n12505_o ? n12512_o : n12565_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12584_o = n12505_o ? n12513_o : n12566_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12585_o = n12505_o ? n12514_o : n12567_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12586_o = n12505_o ? n12515_o : n12568_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12587_o = n12505_o ? n12516_o : n12569_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12588_o = n12505_o ? n12517_o : n12570_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12589_o = n12505_o ? n12506_o : n12571_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12590_o = n12505_o ? n12507_o : n12572_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12591_o = n12505_o ? n12518_o : n12573_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12592_o = n12505_o ? n12519_o : n12574_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12593_o = n12505_o ? n12520_o : n12575_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12594_o = n12505_o ? n12521_o : n12576_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12595_o = n12505_o ? n12522_o : n12577_o;
  /* ../../HW/src/dp/dp_sink.vhd:312:1  */
  assign n12596_o = n12505_o ? n12523_o : n12578_o;
  /* ../../HW/src/dp/dp_sink.vhd:464:17  */
  assign n12638_o = ~reset_in;
  /* ../../HW/src/dp/dp_sink.vhd:515:26  */
  assign n12641_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:515:53  */
  assign n12642_o = wr_datavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:515:34  */
  assign n12643_o = n12642_o & n12641_o;
  /* ../../HW/src/dp/dp_sink.vhd:515:70  */
  assign n12644_o = ~wr_vm;
  /* ../../HW/src/dp/dp_sink.vhd:515:61  */
  assign n12645_o = n12644_o & n12643_o;
  /* ../../HW/src/dp/dp_sink.vhd:516:41  */
  assign n12647_o = req_p0_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:515:13  */
  assign n12648_o = n12645_o ? n12647_o : req_p0_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:520:26  */
  assign n12649_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:520:53  */
  assign n12650_o = wr_datavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:520:34  */
  assign n12651_o = n12650_o & n12649_o;
  /* ../../HW/src/dp/dp_sink.vhd:520:70  */
  assign n12652_o = ~wr_vm;
  /* ../../HW/src/dp/dp_sink.vhd:520:61  */
  assign n12653_o = n12652_o & n12651_o;
  /* ../../HW/src/dp/dp_sink.vhd:521:41  */
  assign n12655_o = req_p0_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:520:13  */
  assign n12656_o = n12653_o ? n12655_o : req_p0_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:525:26  */
  assign n12657_o = wr_req_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:525:53  */
  assign n12658_o = wr_datavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:525:34  */
  assign n12659_o = n12658_o & n12657_o;
  /* ../../HW/src/dp/dp_sink.vhd:525:70  */
  assign n12660_o = ~wr_vm;
  /* ../../HW/src/dp/dp_sink.vhd:525:61  */
  assign n12661_o = n12660_o & n12659_o;
  /* ../../HW/src/dp/dp_sink.vhd:526:41  */
  assign n12663_o = req_p0_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:525:13  */
  assign n12664_o = n12661_o ? n12663_o : req_p0_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:533:26  */
  assign n12665_o = wr_req_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:533:53  */
  assign n12666_o = wr_datavalid_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:533:34  */
  assign n12667_o = n12666_o & n12665_o;
  /* ../../HW/src/dp/dp_sink.vhd:533:61  */
  assign n12668_o = wr_vm & n12667_o;
  /* ../../HW/src/dp/dp_sink.vhd:534:41  */
  assign n12670_o = req_p1_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:533:13  */
  assign n12671_o = n12668_o ? n12670_o : req_p1_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:538:26  */
  assign n12672_o = wr_req_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:538:53  */
  assign n12673_o = wr_datavalid_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:538:34  */
  assign n12674_o = n12673_o & n12672_o;
  /* ../../HW/src/dp/dp_sink.vhd:538:61  */
  assign n12675_o = wr_vm & n12674_o;
  /* ../../HW/src/dp/dp_sink.vhd:539:41  */
  assign n12677_o = req_p1_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:538:13  */
  assign n12678_o = n12675_o ? n12677_o : req_p1_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:543:26  */
  assign n12679_o = wr_req_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:543:53  */
  assign n12680_o = wr_datavalid_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:543:34  */
  assign n12681_o = n12680_o & n12679_o;
  /* ../../HW/src/dp/dp_sink.vhd:543:61  */
  assign n12682_o = wr_vm & n12681_o;
  /* ../../HW/src/dp/dp_sink.vhd:544:41  */
  assign n12684_o = req_p1_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:543:13  */
  assign n12685_o = n12682_o ? n12684_o : req_p1_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:551:23  */
  assign n12686_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:551:57  */
  assign n12687_o = wr_readdatavalid_vm_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:551:60  */
  assign n12688_o = ~n12687_o;
  /* ../../HW/src/dp/dp_sink.vhd:551:31  */
  assign n12689_o = n12688_o & n12686_o;
  /* ../../HW/src/dp/dp_sink.vhd:552:41  */
  assign n12691_o = rsp_p0_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:551:13  */
  assign n12692_o = n12689_o ? n12691_o : rsp_p0_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:556:23  */
  assign n12693_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:556:57  */
  assign n12694_o = wr_readdatavalid_vm_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:556:60  */
  assign n12695_o = ~n12694_o;
  /* ../../HW/src/dp/dp_sink.vhd:556:31  */
  assign n12696_o = n12695_o & n12693_o;
  /* ../../HW/src/dp/dp_sink.vhd:557:41  */
  assign n12698_o = rsp_p0_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:556:13  */
  assign n12699_o = n12696_o ? n12698_o : rsp_p0_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:561:23  */
  assign n12700_o = wr_req2[2];
  /* ../../HW/src/dp/dp_sink.vhd:561:57  */
  assign n12701_o = wr_readdatavalid_vm_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:561:60  */
  assign n12702_o = ~n12701_o;
  /* ../../HW/src/dp/dp_sink.vhd:561:31  */
  assign n12703_o = n12702_o & n12700_o;
  /* ../../HW/src/dp/dp_sink.vhd:562:41  */
  assign n12705_o = rsp_p0_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:561:13  */
  assign n12706_o = n12703_o ? n12705_o : rsp_p0_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:569:23  */
  assign n12707_o = wr_req2[0];
  /* ../../HW/src/dp/dp_sink.vhd:569:57  */
  assign n12708_o = wr_readdatavalid_vm_in[0];
  /* ../../HW/src/dp/dp_sink.vhd:569:31  */
  assign n12709_o = n12708_o & n12707_o;
  /* ../../HW/src/dp/dp_sink.vhd:570:41  */
  assign n12711_o = rsp_p1_0_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:569:13  */
  assign n12712_o = n12709_o ? n12711_o : rsp_p1_0_r;
  /* ../../HW/src/dp/dp_sink.vhd:574:23  */
  assign n12713_o = wr_req2[1];
  /* ../../HW/src/dp/dp_sink.vhd:574:57  */
  assign n12714_o = wr_readdatavalid_vm_in[1];
  /* ../../HW/src/dp/dp_sink.vhd:574:31  */
  assign n12715_o = n12714_o & n12713_o;
  /* ../../HW/src/dp/dp_sink.vhd:575:41  */
  assign n12717_o = rsp_p1_1_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:574:13  */
  assign n12718_o = n12715_o ? n12717_o : rsp_p1_1_r;
  /* ../../HW/src/dp/dp_sink.vhd:579:23  */
  assign n12719_o = wr_req2[2];
  /* ../../HW/src/dp/dp_sink.vhd:579:57  */
  assign n12720_o = wr_readdatavalid_vm_in[2];
  /* ../../HW/src/dp/dp_sink.vhd:579:31  */
  assign n12721_o = n12720_o & n12719_o;
  /* ../../HW/src/dp/dp_sink.vhd:580:41  */
  assign n12723_o = rsp_p1_2_r + 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:579:13  */
  assign n12724_o = n12721_o ? n12723_o : rsp_p1_2_r;
  /* ../../HW/src/dp/dp_sink.vhd:601:28  */
  assign n12725_o = n12648_o != n12692_o;
  /* ../../HW/src/dp/dp_sink.vhd:601:13  */
  assign n12728_o = n12725_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:607:28  */
  assign n12729_o = n12656_o != n12699_o;
  /* ../../HW/src/dp/dp_sink.vhd:607:13  */
  assign n12732_o = n12729_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:613:28  */
  assign n12733_o = n12664_o != n12706_o;
  /* ../../HW/src/dp/dp_sink.vhd:613:13  */
  assign n12736_o = n12733_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:621:28  */
  assign n12737_o = n12671_o != n12712_o;
  /* ../../HW/src/dp/dp_sink.vhd:621:13  */
  assign n12740_o = n12737_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:627:28  */
  assign n12741_o = n12678_o != n12718_o;
  /* ../../HW/src/dp/dp_sink.vhd:627:13  */
  assign n12744_o = n12741_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:633:28  */
  assign n12745_o = n12685_o != n12724_o;
  /* ../../HW/src/dp/dp_sink.vhd:633:13  */
  assign n12748_o = n12745_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:639:35  */
  assign n12749_o = ~bus_wait_request_in;
  /* ../../HW/src/dp/dp_sink.vhd:639:51  */
  assign n12750_o = ~valid_rr;
  /* ../../HW/src/dp/dp_sink.vhd:639:40  */
  assign n12751_o = n12749_o | n12750_o;
  /* ../../HW/src/dp/dp_sink.vhd:647:23  */
  assign n12752_o = q_r[0];
  /* ../../HW/src/dp/dp_sink.vhd:651:98  */
  assign n12753_o = q_r[64:1];
  /* ../../HW/src/dp/dp_sink.vhd:647:17  */
  assign n12754_o = n12752_o ? q2 : n12753_o;
  /* ../../HW/src/dp/dp_sink.vhd:656:49  */
  assign n12755_o = q_r[96:65];
  /* ../../HW/src/dp/dp_sink.vhd:659:34  */
  assign n12756_o = q_r[97];
  /* ../../HW/src/dp/dp_sink.vhd:661:39  */
  assign n12757_o = q_r[98];
  /* ../../HW/src/dp/dp_sink.vhd:663:32  */
  assign n12758_o = q_r[99];
  /* ../../HW/src/dp/dp_sink.vhd:681:41  */
  assign n12759_o = q_r[106:105];
  /* ../../HW/src/dp/dp_sink.vhd:683:45  */
  assign n12760_o = q_r[107];
  /* ../../HW/src/dp/dp_sink.vhd:685:48  */
  assign n12761_o = q_r[109:108];
  /* ../../HW/src/dp/dp_sink.vhd:687:40  */
  assign n12762_o = q_r[111:110];
  /* ../../HW/src/dp/dp_sink.vhd:689:52  */
  assign n12763_o = q_r[117:112];
  /* ../../HW/src/dp/dp_sink.vhd:691:32  */
  assign n12764_o = q_r[120:118];
  /* ../../HW/src/dp/dp_sink.vhd:693:32  */
  assign n12765_o = q_r[121];
  /* ../../HW/src/dp/dp_sink.vhd:695:44  */
  assign n12766_o = q_r[123:122];
  /* ../../HW/src/dp/dp_sink.vhd:697:33  */
  assign n12767_o = q_r[125:124];
  /* ../../HW/src/dp/dp_sink.vhd:699:35  */
  assign n12768_o = q_r[127:126];
  /* ../../HW/src/dp/dp_sink.vhd:702:44  */
  assign n12769_o = q_r[131:128];
  /* ../../HW/src/dp/dp_sink.vhd:706:38  */
  assign n12773_o = n12764_o == 3'b001;
  /* ../../HW/src/dp/dp_sink.vhd:707:35  */
  assign n12775_o = $unsigned(9'b000000001) > $unsigned(9'b000010100);
  /* ../../HW/src/dp/dp_sink.vhd:707:20  */
  assign n12777_o = n12775_o ? 9'b000010011 : 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:710:50  */
  assign n12778_o = n12777_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:711:51  */
  assign n12780_o = n12777_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_sink.vhd:712:41  */
  assign n12782_o = n12764_o == 3'b011;
  /* ../../HW/src/dp/dp_sink.vhd:713:35  */
  assign n12784_o = $unsigned(9'b000000001) > $unsigned(9'b000001010);
  /* ../../HW/src/dp/dp_sink.vhd:713:20  */
  assign n12786_o = n12784_o ? 9'b000001001 : 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:716:50  */
  assign n12787_o = n12786_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:717:51  */
  assign n12789_o = n12786_o << 32'b00000000000000000000000000000010;
  /* ../../HW/src/dp/dp_sink.vhd:718:41  */
  assign n12791_o = n12764_o == 3'b111;
  /* ../../HW/src/dp/dp_sink.vhd:719:35  */
  assign n12793_o = $unsigned(9'b000000001) > $unsigned(9'b000000101);
  /* ../../HW/src/dp/dp_sink.vhd:719:20  */
  assign n12795_o = n12793_o ? 9'b000000100 : 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:722:50  */
  assign n12796_o = n12795_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:723:51  */
  assign n12798_o = n12795_o << 32'b00000000000000000000000000000011;
  /* ../../HW/src/dp/dp_sink.vhd:725:35  */
  assign n12800_o = $unsigned(9'b000000001) > $unsigned(9'b000101000);
  /* ../../HW/src/dp/dp_sink.vhd:725:20  */
  assign n12802_o = n12800_o ? 9'b000100111 : 9'b000000001;
  /* ../../HW/src/dp/dp_sink.vhd:728:50  */
  assign n12803_o = n12802_o[4:0];
  /* ../../HW/src/dp/dp_sink.vhd:718:17  */
  assign n12804_o = n12791_o ? n12798_o : n12802_o;
  /* ../../HW/src/dp/dp_sink.vhd:718:17  */
  assign n12805_o = n12791_o ? n12796_o : n12803_o;
  /* ../../HW/src/dp/dp_sink.vhd:712:17  */
  assign n12807_o = n12782_o ? n12789_o : n12804_o;
  /* ../../HW/src/dp/dp_sink.vhd:712:17  */
  assign n12808_o = n12782_o ? n12787_o : n12805_o;
  /* ../../HW/src/dp/dp_sink.vhd:706:17  */
  assign n12810_o = n12773_o ? n12780_o : n12807_o;
  /* ../../HW/src/dp/dp_sink.vhd:706:17  */
  assign n12811_o = n12773_o ? n12778_o : n12808_o;
  assign n12890_o = {n12736_o, n12732_o, n12728_o};
  assign n12892_o = {n12748_o, n12744_o, n12740_o};
  /* ../../HW/src/dp/dp_sink.vhd:759:12  */
  assign n13151_o = ~reset_in;
  /* ../../HW/src/dp/dp_sink.vhd:764:27  */
  assign n13153_o = ~usedw;
  /* ../../HW/src/dp/dp_sink.vhd:765:18  */
  assign n13155_o = $unsigned(n13153_o) <= $unsigned(9'b000101111);
  /* ../../HW/src/dp/dp_sink.vhd:765:7  */
  assign n13158_o = n13155_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:775:26  */
  assign n13173_o = ~empty;
  /* ../../HW/src/dp/dp_sink.vhd:775:44  */
  assign n13174_o = ~empty2;
  /* ../../HW/src/dp/dp_sink.vhd:775:54  */
  assign n13175_o = q[0];
  /* ../../HW/src/dp/dp_sink.vhd:775:57  */
  assign n13176_o = ~n13175_o;
  /* ../../HW/src/dp/dp_sink.vhd:775:50  */
  assign n13177_o = n13174_o | n13176_o;
  /* ../../HW/src/dp/dp_sink.vhd:775:32  */
  assign n13178_o = n13177_o & n13173_o;
  /* ../../HW/src/dp/dp_sink.vhd:775:15  */
  assign n13179_o = n13178_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:787:20  */
  assign n13183_o = q[0];
  /* ../../HW/src/dp/dp_sink.vhd:784:5  */
  assign n13185_o = emptyn ? emptyn : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:784:5  */
  assign n13187_o = emptyn ? n13183_o : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:784:5  */
  assign n13190_o = emptyn ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:780:5  */
  assign n13192_o = bus_wait_request_in ? 1'b0 : n13185_o;
  /* ../../HW/src/dp/dp_sink.vhd:780:5  */
  assign n13194_o = bus_wait_request_in ? 1'b0 : n13187_o;
  /* ../../HW/src/dp/dp_sink.vhd:780:5  */
  assign n13195_o = bus_wait_request_in ? valid_r : n13190_o;
  /* ../../HW/src/dp/dp_sink.vhd:797:20  */
  assign n13196_o = q[0];
  /* ../../HW/src/dp/dp_sink.vhd:794:5  */
  assign n13198_o = emptyn ? emptyn : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:794:5  */
  assign n13200_o = emptyn ? n13196_o : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:794:5  */
  assign n13203_o = emptyn ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_sink.vhd:779:1  */
  assign n13204_o = valid_rr ? n13192_o : n13198_o;
  /* ../../HW/src/dp/dp_sink.vhd:779:1  */
  assign n13205_o = valid_rr ? n13194_o : n13200_o;
  /* ../../HW/src/dp/dp_sink.vhd:779:1  */
  assign n13206_o = valid_rr ? n13195_o : n13203_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13210_o = rdreq ? q : q_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13211_q <= 132'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n13211_q <= n13210_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13212_o = n12751_o ? valid : valid_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13213_q <= 1'b0;
    else
      n13213_q <= n13212_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13214_o = n12751_o ? valid_r : valid_rr;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13215_q <= 1'b0;
    else
      n13215_q <= n13214_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13216_o = n12751_o ? n12768_o : bus_data_flow_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13217_q <= 2'b00;
    else
      n13217_q <= n13216_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13218_o = n12751_o ? n12769_o : bus_end_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13219_q <= 4'b0000;
    else
      n13219_q <= n13218_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13220_o = n12751_o ? n12764_o : bus_vector_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13221_q <= 3'b000;
    else
      n13221_q <= n13220_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13222_o = n12751_o ? n12765_o : bus_stream_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13223_q <= 1'b0;
    else
      n13223_q <= n13222_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13224_o = n12751_o ? n12766_o : bus_stream_id_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13225_q <= 2'b00;
    else
      n13225_q <= n13224_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13226_o = n12751_o ? n12767_o : bus_scatter_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13227_q <= 2'b00;
    else
      n13227_q <= n13226_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13228_o = n12751_o ? n12755_o : bus_addr_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13229_q <= 32'b00000000000000000000000000000000;
    else
      n13229_q <= n13228_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13230_o = n12751_o ? n12756_o : bus_fork_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13231_q <= 1'b0;
    else
      n13231_q <= n13230_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13232_o = n12751_o ? n12757_o : bus_addr_mode_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13233_q <= 1'b0;
    else
      n13233_q <= n13232_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13234_o = n12751_o ? n12758_o : bus_vm_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13235_q <= 1'b0;
    else
      n13235_q <= n13234_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13236_o = n12751_o ? n12754_o : bus_writedata_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13237_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n13237_q <= n13236_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13238_o = n12751_o ? 5'b00001 : bus_burstlen_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13239_q <= 5'b00000;
    else
      n13239_q <= n13238_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13240_o = n12751_o ? n12810_o : bus_burstlen2_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13241_q <= 9'b000000000;
    else
      n13241_q <= n13240_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13242_o = n12751_o ? n12811_o : bus_burstlen3_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13243_q <= 5'b00000;
    else
      n13243_q <= n13242_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13244_o = n12751_o ? n12759_o : bus_id_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13245_q <= 2'b00;
    else
      n13245_q <= n13244_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13246_o = n12751_o ? n12760_o : bus_thread_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13247_q <= 1'b0;
    else
      n13247_q <= n13246_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13248_o = n12751_o ? n12761_o : bus_data_type_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13249_q <= 2'b00;
    else
      n13249_q <= n13248_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13250_o = n12751_o ? n12762_o : bus_data_model_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13251_q <= 2'b00;
    else
      n13251_q <= n13250_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  assign n13252_o = n12751_o ? n12763_o : bus_mcast_r;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13253_q <= 6'b111111;
    else
      n13253_q <= n13252_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13254_q <= 9'b000000000;
    else
      n13254_q <= n12648_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13255_q <= 9'b000000000;
    else
      n13255_q <= n12656_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13256_q <= 9'b000000000;
    else
      n13256_q <= n12664_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13257_q <= 9'b000000000;
    else
      n13257_q <= n12692_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13258_q <= 9'b000000000;
    else
      n13258_q <= n12699_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13259_q <= 9'b000000000;
    else
      n13259_q <= n12706_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13260_q <= 9'b000000000;
    else
      n13260_q <= n12671_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13261_q <= 9'b000000000;
    else
      n13261_q <= n12678_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13262_q <= 9'b000000000;
    else
      n13262_q <= n12685_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13263_q <= 9'b000000000;
    else
      n13263_q <= n12712_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13264_q <= 9'b000000000;
    else
      n13264_q <= n12718_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13265_q <= 9'b000000000;
    else
      n13265_q <= n12724_o;
  /* ../../HW/src/dp/dp_sink.vhd:464:5  */
  assign n13266_o = {wr_end, wr_data_flow, wr_scatter, wr_stream_id, wr_stream, wr_vector, wr_mcast, wr_data_model, wr_data_type, wr_thread, wr_bus_id, wr_burstlen, wr_vm, wr_addr_mode, wr_fork, wr_addr, wr_data, wr_datavalid};
  /* ../../HW/src/dp/dp_sink.vhd:464:5  */
  assign n13267_o = {n12484_o, n12476_o, n12468_o};
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13268_q <= 3'b000;
    else
      n13268_q <= n12890_o;
  /* ../../HW/src/dp/dp_sink.vhd:504:9  */
  always @(posedge clock_in or posedge n12638_o)
    if (n12638_o)
      n13269_q <= 3'b000;
    else
      n13269_q <= n12892_o;
  /* ../../HW/src/dp/dp_sink.vhd:763:4  */
  always @(posedge clock_in or posedge n13151_o)
    if (n13151_o)
      n13270_q <= 1'b0;
    else
      n13270_q <= n13158_o;
  /* ../../HW/src/dp/dp_sink.vhd:763:4  */
  always @(posedge clock_in or posedge n13151_o)
    if (n13151_o)
      n13271_q <= 5'b00000;
    else
      n13271_q <= 5'b11111;
endmodule

module dp_source_2_3_1_32_1_0
  (input  clock_in,
   input  reset_in,
   input  bus_readdatavalid_in,
   input  bus_readdatavalid_vm_in,
   input  [63:0] bus_readdata_in,
   input  bus_wait_request_in,
   input  gen_valid_in,
   input  gen_vm_in,
   input  gen_fork_in,
   input  [1:0] gen_data_flow_in,
   input  gen_src_stream_in,
   input  gen_dest_stream_in,
   input  [1:0] gen_stream_id_in,
   input  [2:0] gen_src_vector_in,
   input  [2:0] gen_dst_vector_in,
   input  [1:0] gen_src_scatter_in,
   input  [1:0] gen_dst_scatter_in,
   input  [3:0] gen_src_start_in,
   input  [3:0] gen_src_end_in,
   input  [3:0] gen_dst_end_in,
   input  gen_src_eof_in,
   input  [31:0] gen_src_addr_in,
   input  gen_src_addr_mode_in,
   input  [31:0] gen_dst_addr_in,
   input  gen_dst_addr_mode_in,
   input  [1:0] gen_bus_id_source_in,
   input  [1:0] gen_data_type_source_in,
   input  [1:0] gen_data_model_source_in,
   input  [1:0] gen_bus_id_dest_in,
   input  gen_busy_dest_in,
   input  [1:0] gen_data_type_dest_in,
   input  [1:0] gen_data_model_dest_in,
   input  [4:0] gen_src_burstlen_in,
   input  [4:0] gen_dst_burstlen_in,
   input  gen_thread_in,
   input  [5:0] gen_mcast_in,
   input  [63:0] gen_src_data_in,
   input  [2:0] wr_full_in,
   output [31:0] bus_addr_out,
   output bus_addr_mode_out,
   output bus_cs_out,
   output bus_read_out,
   output bus_read_vm_out,
   output bus_read_fork_out,
   output [1:0] bus_read_data_flow_out,
   output bus_read_stream_out,
   output [1:0] bus_read_stream_id_out,
   output [2:0] bus_read_vector_out,
   output [1:0] bus_read_scatter_out,
   output [3:0] bus_read_start_out,
   output [3:0] bus_read_end_out,
   output [4:0] bus_burstlen_out,
   output [1:0] bus_id_out,
   output [1:0] bus_data_type_out,
   output [1:0] bus_data_model_out,
   output gen_waitreq_out,
   output [2:0] wr_req_out,
   output [2:0] wr_req_pending_p0_out,
   output [2:0] wr_req_pending_p1_out,
   output [5:0] wr_data_flow_out,
   output [8:0] wr_vector_out,
   output [2:0] wr_stream_out,
   output [5:0] wr_stream_id_out,
   output [5:0] wr_scatter_out,
   output [11:0] wr_end_out,
   output [31:0] wr_addr_out,
   output wr_fork_out,
   output wr_addr_mode_out,
   output wr_src_vm_out,
   output wr_datavalid_out,
   output [63:0] wr_data_out,
   output wr_readdatavalid_out,
   output wr_readdatavalid_vm_out,
   output [63:0] wr_readdata_out,
   output [4:0] wr_burstlen_out,
   output [1:0] wr_bus_id_out,
   output wr_thread_out,
   output [1:0] wr_data_type_out,
   output [1:0] wr_data_model_out,
   output [5:0] wr_mcast_out);
  wire doit;
  wire wr_req;
  wire [31:0] wr_addr;
  wire wr_fork;
  wire wr_addr_mode;
  wire wr_src_vm;
  wire [1:0] dp_bus_id;
  wire [1:0] dp_data_type;
  wire [1:0] dp_data_model;
  wire dp_thread;
  wire [5:0] dp_mcast;
  wire [4:0] wr_burstlen;
  wire gen_valid;
  wire [63:0] bus_readdata;
  wire n12259_o;
  wire n12260_o;
  wire [63:0] n12261_o;
  localparam n12264_o = 1'b1;
  wire delay_i1_out_out;
  localparam n12268_o = 1'b1;
  wire [1:0] delay_i3_out_out;
  localparam n12272_o = 1'b1;
  wire [1:0] delay_i4_out_out;
  localparam n12276_o = 1'b1;
  wire delay_i5_out_out;
  localparam n12280_o = 1'b1;
  wire [4:0] delay_i6_out_out;
  localparam n12284_o = 1'b1;
  wire [5:0] delay_i7_out_out;
  localparam n12288_o = 1'b1;
  wire delay_i8_out_out;
  localparam n12292_o = 1'b1;
  wire [63:0] delay_i9_out_out;
  localparam n12296_o = 1'b1;
  wire [63:0] gen_delay_i10_out_out;
  wire n12300_o;
  wire n12301_o;
  wire n12302_o;
  wire n12303_o;
  wire n12304_o;
  wire n12305_o;
  wire n12306_o;
  wire n12308_o;
  wire n12309_o;
  wire n12310_o;
  wire n12311_o;
  wire n12314_o;
  wire [30:0] n12317_o;
  wire [31:0] n12318_o;
  wire n12320_o;
  wire n12322_o;
  wire [30:0] n12323_o;
  wire [31:0] n12324_o;
  wire n12326_o;
  wire n12327_o;
  wire n12328_o;
  wire n12330_o;
  wire [30:0] n12331_o;
  wire [31:0] n12332_o;
  wire n12334_o;
  wire n12335_o;
  wire n12337_o;
  wire [30:0] n12338_o;
  wire [31:0] n12339_o;
  wire n12341_o;
  wire n12343_o;
  wire [30:0] n12344_o;
  wire [31:0] n12345_o;
  wire n12347_o;
  wire n12348_o;
  wire n12349_o;
  wire n12351_o;
  wire [30:0] n12352_o;
  wire [31:0] n12353_o;
  wire n12355_o;
  wire n12356_o;
  wire n12358_o;
  wire [30:0] n12359_o;
  wire [31:0] n12360_o;
  wire n12362_o;
  wire n12364_o;
  wire [30:0] n12365_o;
  wire [31:0] n12366_o;
  wire n12368_o;
  wire n12369_o;
  wire n12370_o;
  wire n12372_o;
  wire [30:0] n12373_o;
  wire [31:0] n12374_o;
  wire n12376_o;
  wire n12377_o;
  wire n12379_o;
  wire n12383_o;
  wire n12384_o;
  wire n12385_o;
  wire n12388_o;
  wire [2:0] n12390_o;
  wire [2:0] n12391_o;
  wire [2:0] n12392_o;
  wire [5:0] n12393_o;
  wire [8:0] n12394_o;
  wire [2:0] n12395_o;
  wire [5:0] n12396_o;
  wire [5:0] n12397_o;
  wire [11:0] n12398_o;
  assign bus_addr_out = gen_src_addr_in;
  assign bus_addr_mode_out = gen_src_addr_mode_in;
  assign bus_cs_out = n12309_o;
  assign bus_read_out = n12311_o;
  assign bus_read_vm_out = gen_vm_in;
  assign bus_read_fork_out = gen_fork_in;
  assign bus_read_data_flow_out = gen_data_flow_in;
  assign bus_read_stream_out = gen_src_stream_in;
  assign bus_read_stream_id_out = gen_stream_id_in;
  assign bus_read_vector_out = gen_src_vector_in;
  assign bus_read_scatter_out = gen_src_scatter_in;
  assign bus_read_start_out = gen_src_start_in;
  assign bus_read_end_out = gen_src_end_in;
  assign bus_burstlen_out = gen_src_burstlen_in;
  assign bus_id_out = gen_bus_id_source_in;
  assign bus_data_type_out = gen_data_type_source_in;
  assign bus_data_model_out = gen_data_model_source_in;
  assign gen_waitreq_out = n12306_o;
  assign wr_req_out = n12390_o;
  assign wr_req_pending_p0_out = n12391_o;
  assign wr_req_pending_p1_out = n12392_o;
  assign wr_data_flow_out = n12393_o;
  assign wr_vector_out = n12394_o;
  assign wr_stream_out = n12395_o;
  assign wr_stream_id_out = n12396_o;
  assign wr_scatter_out = n12397_o;
  assign wr_end_out = n12398_o;
  assign wr_addr_out = wr_addr;
  assign wr_fork_out = wr_fork;
  assign wr_addr_mode_out = wr_addr_mode;
  assign wr_src_vm_out = wr_src_vm;
  assign wr_datavalid_out = n12314_o;
  assign wr_data_out = gen_src_data_in;
  assign wr_readdatavalid_out = bus_readdatavalid_in;
  assign wr_readdatavalid_vm_out = bus_readdatavalid_vm_in;
  assign wr_readdata_out = bus_readdata;
  assign wr_burstlen_out = wr_burstlen;
  assign wr_bus_id_out = dp_bus_id;
  assign wr_thread_out = dp_thread;
  assign wr_data_type_out = dp_data_type;
  assign wr_data_model_out = dp_data_model;
  assign wr_mcast_out = dp_mcast;
  /* ../../HW/src/dp/dp_source.vhd:135:8  */
  assign doit = gen_valid; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:136:8  */
  assign wr_req = n12388_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:137:8  */
  assign wr_addr = gen_dst_addr_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:138:8  */
  assign wr_fork = gen_fork_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:139:8  */
  assign wr_addr_mode = gen_dst_addr_mode_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:140:8  */
  assign wr_src_vm = gen_vm_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:141:8  */
  assign dp_bus_id = gen_bus_id_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:142:8  */
  assign dp_data_type = gen_data_type_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:143:8  */
  assign dp_data_model = gen_data_model_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:144:8  */
  assign dp_thread = gen_thread_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:145:8  */
  assign dp_mcast = gen_mcast_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:146:8  */
  assign wr_burstlen = gen_dst_burstlen_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:155:8  */
  assign gen_valid = n12260_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:156:8  */
  assign bus_readdata = n12261_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:160:32  */
  assign n12259_o = ~gen_busy_dest_in;
  /* ../../HW/src/dp/dp_source.vhd:160:27  */
  assign n12260_o = gen_valid_in & n12259_o;
  /* ../../HW/src/dp/dp_source.vhd:162:33  */
  assign n12261_o = bus_readdatavalid_in ? bus_readdata_in : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/dp/dp_source.vhd:164:1  */
  delay_8 delay_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_req),
    .enable_in(n12264_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:166:1  */
  delayi_2_8 delay_i3 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_bus_id),
    .enable_in(n12268_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:168:1  */
  delayi_2_8 delay_i4 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_data_type),
    .enable_in(n12272_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:170:1  */
  delayi_1_8 delay_i5 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_thread),
    .enable_in(n12276_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:172:1  */
  delayi_5_8 delay_i6 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_burstlen),
    .enable_in(n12280_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:174:1  */
  delayv_6_8 delay_i7 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_mcast),
    .enable_in(n12284_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:176:1  */
  delay_8 delay_i8 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(gen_src_eof_in),
    .enable_in(n12288_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:178:1  */
  delayv_64_8 delay_i9 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(gen_src_data_in),
    .enable_in(n12292_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:182:1  */
  delayv_64_7 gen_delay_i10 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(bus_readdata),
    .enable_in(n12296_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:190:39  */
  assign n12300_o = bus_wait_request_in & doit;
  /* ../../HW/src/dp/dp_source.vhd:190:85  */
  assign n12301_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:190:67  */
  assign n12302_o = n12301_o & n12300_o;
  /* ../../HW/src/dp/dp_source.vhd:190:104  */
  assign n12303_o = ~gen_valid;
  /* ../../HW/src/dp/dp_source.vhd:190:109  */
  assign n12304_o = gen_valid_in & n12303_o;
  /* ../../HW/src/dp/dp_source.vhd:190:91  */
  assign n12305_o = n12302_o | n12304_o;
  /* ../../HW/src/dp/dp_source.vhd:190:24  */
  assign n12306_o = n12305_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:202:30  */
  assign n12308_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:202:25  */
  assign n12309_o = gen_valid & n12308_o;
  /* ../../HW/src/dp/dp_source.vhd:203:32  */
  assign n12310_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:203:27  */
  assign n12311_o = gen_valid & n12310_o;
  /* ../../HW/src/dp/dp_source.vhd:234:21  */
  assign n12314_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n12317_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12318_o = {1'b0, n12317_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12320_o = 32'b00000000000000000000000000000000 == n12318_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12322_o = n12320_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12323_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12324_o = {1'b0, n12323_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12326_o = 32'b00000000000000000000000000000000 == n12324_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12327_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12328_o = gen_valid_in & n12327_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12330_o = n12326_o ? n12328_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12331_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12332_o = {1'b0, n12331_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12334_o = 32'b00000000000000000000000000000000 == n12332_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12335_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12337_o = n12334_o ? n12335_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n12338_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12339_o = {1'b0, n12338_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12341_o = 32'b00000000000000000000000000000001 == n12339_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12343_o = n12341_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12344_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12345_o = {1'b0, n12344_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12347_o = 32'b00000000000000000000000000000001 == n12345_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12348_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12349_o = gen_valid_in & n12348_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12351_o = n12347_o ? n12349_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12352_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12353_o = {1'b0, n12352_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12355_o = 32'b00000000000000000000000000000001 == n12353_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12356_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12358_o = n12355_o ? n12356_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n12359_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12360_o = {1'b0, n12359_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12362_o = 32'b00000000000000000000000000000010 == n12360_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12364_o = n12362_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12365_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12366_o = {1'b0, n12365_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12368_o = 32'b00000000000000000000000000000010 == n12366_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12369_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12370_o = gen_valid_in & n12369_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12372_o = n12368_o ? n12370_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12373_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12374_o = {1'b0, n12373_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12376_o = 32'b00000000000000000000000000000010 == n12374_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12377_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12379_o = n12376_o ? n12377_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:278:41  */
  assign n12383_o = ~bus_wait_request_in;
  /* ../../HW/src/dp/dp_source.vhd:278:46  */
  assign n12384_o = n12383_o | gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:278:17  */
  assign n12385_o = n12384_o & doit;
  /* ../../HW/src/dp/dp_source.vhd:278:5  */
  assign n12388_o = n12385_o ? 1'b1 : 1'b0;
  assign n12390_o = {n12364_o, n12343_o, n12322_o};
  assign n12391_o = {n12372_o, n12351_o, n12330_o};
  assign n12392_o = {n12379_o, n12358_o, n12337_o};
  assign n12393_o = {gen_data_flow_in, gen_data_flow_in, gen_data_flow_in};
  assign n12394_o = {gen_dst_vector_in, gen_dst_vector_in, gen_dst_vector_in};
  assign n12395_o = {gen_dest_stream_in, gen_dest_stream_in, gen_dest_stream_in};
  assign n12396_o = {gen_stream_id_in, gen_stream_id_in, gen_stream_id_in};
  assign n12397_o = {gen_dst_scatter_in, gen_dst_scatter_in, gen_dst_scatter_in};
  assign n12398_o = {gen_dst_end_in, gen_dst_end_in, gen_dst_end_in};
endmodule

module dp_source_1_3_4_32_1_0
  (input  clock_in,
   input  reset_in,
   input  bus_readdatavalid_in,
   input  bus_readdatavalid_vm_in,
   input  [63:0] bus_readdata_in,
   input  bus_wait_request_in,
   input  gen_valid_in,
   input  gen_vm_in,
   input  gen_fork_in,
   input  [1:0] gen_data_flow_in,
   input  gen_src_stream_in,
   input  gen_dest_stream_in,
   input  [1:0] gen_stream_id_in,
   input  [2:0] gen_src_vector_in,
   input  [2:0] gen_dst_vector_in,
   input  [1:0] gen_src_scatter_in,
   input  [1:0] gen_dst_scatter_in,
   input  [3:0] gen_src_start_in,
   input  [3:0] gen_src_end_in,
   input  [3:0] gen_dst_end_in,
   input  gen_src_eof_in,
   input  [31:0] gen_src_addr_in,
   input  gen_src_addr_mode_in,
   input  [31:0] gen_dst_addr_in,
   input  gen_dst_addr_mode_in,
   input  [1:0] gen_bus_id_source_in,
   input  [1:0] gen_data_type_source_in,
   input  [1:0] gen_data_model_source_in,
   input  [1:0] gen_bus_id_dest_in,
   input  gen_busy_dest_in,
   input  [1:0] gen_data_type_dest_in,
   input  [1:0] gen_data_model_dest_in,
   input  [4:0] gen_src_burstlen_in,
   input  [4:0] gen_dst_burstlen_in,
   input  gen_thread_in,
   input  [5:0] gen_mcast_in,
   input  [63:0] gen_src_data_in,
   input  [2:0] wr_full_in,
   output [31:0] bus_addr_out,
   output bus_addr_mode_out,
   output bus_cs_out,
   output bus_read_out,
   output bus_read_vm_out,
   output bus_read_fork_out,
   output [1:0] bus_read_data_flow_out,
   output bus_read_stream_out,
   output [1:0] bus_read_stream_id_out,
   output [2:0] bus_read_vector_out,
   output [1:0] bus_read_scatter_out,
   output [3:0] bus_read_start_out,
   output [3:0] bus_read_end_out,
   output [4:0] bus_burstlen_out,
   output [1:0] bus_id_out,
   output [1:0] bus_data_type_out,
   output [1:0] bus_data_model_out,
   output gen_waitreq_out,
   output [2:0] wr_req_out,
   output [2:0] wr_req_pending_p0_out,
   output [2:0] wr_req_pending_p1_out,
   output [5:0] wr_data_flow_out,
   output [8:0] wr_vector_out,
   output [2:0] wr_stream_out,
   output [5:0] wr_stream_id_out,
   output [5:0] wr_scatter_out,
   output [11:0] wr_end_out,
   output [31:0] wr_addr_out,
   output wr_fork_out,
   output wr_addr_mode_out,
   output wr_src_vm_out,
   output wr_datavalid_out,
   output [63:0] wr_data_out,
   output wr_readdatavalid_out,
   output wr_readdatavalid_vm_out,
   output [63:0] wr_readdata_out,
   output [4:0] wr_burstlen_out,
   output [1:0] wr_bus_id_out,
   output wr_thread_out,
   output [1:0] wr_data_type_out,
   output [1:0] wr_data_model_out,
   output [5:0] wr_mcast_out);
  wire doit;
  wire wr_req;
  wire [31:0] wr_addr;
  wire wr_fork;
  wire wr_addr_mode;
  wire wr_src_vm;
  wire [1:0] dp_bus_id;
  wire [1:0] dp_data_type;
  wire [1:0] dp_data_model;
  wire dp_thread;
  wire [5:0] dp_mcast;
  wire [4:0] wr_burstlen;
  wire gen_valid;
  wire [63:0] bus_readdata;
  wire n12077_o;
  wire n12078_o;
  wire [63:0] n12079_o;
  localparam n12082_o = 1'b1;
  wire delay_i1_out_out;
  localparam n12086_o = 1'b1;
  wire [1:0] delay_i3_out_out;
  localparam n12090_o = 1'b1;
  wire [1:0] delay_i4_out_out;
  localparam n12094_o = 1'b1;
  wire delay_i5_out_out;
  localparam n12098_o = 1'b1;
  wire [4:0] delay_i6_out_out;
  localparam n12102_o = 1'b1;
  wire [5:0] delay_i7_out_out;
  localparam n12106_o = 1'b1;
  wire delay_i8_out_out;
  localparam n12110_o = 1'b1;
  wire [63:0] delay_i9_out_out;
  localparam n12114_o = 1'b1;
  wire [63:0] gen_delay_i10_out_out;
  wire n12118_o;
  wire n12119_o;
  wire n12120_o;
  wire n12121_o;
  wire n12122_o;
  wire n12123_o;
  wire n12124_o;
  wire n12126_o;
  wire n12127_o;
  wire n12128_o;
  wire n12129_o;
  wire n12132_o;
  wire [30:0] n12135_o;
  wire [31:0] n12136_o;
  wire n12138_o;
  wire n12140_o;
  wire [30:0] n12141_o;
  wire [31:0] n12142_o;
  wire n12144_o;
  wire n12145_o;
  wire n12146_o;
  wire n12148_o;
  wire [30:0] n12149_o;
  wire [31:0] n12150_o;
  wire n12152_o;
  wire n12153_o;
  wire n12155_o;
  wire [30:0] n12156_o;
  wire [31:0] n12157_o;
  wire n12159_o;
  wire n12161_o;
  wire [30:0] n12162_o;
  wire [31:0] n12163_o;
  wire n12165_o;
  wire n12166_o;
  wire n12167_o;
  wire n12169_o;
  wire [30:0] n12170_o;
  wire [31:0] n12171_o;
  wire n12173_o;
  wire n12174_o;
  wire n12176_o;
  wire [30:0] n12177_o;
  wire [31:0] n12178_o;
  wire n12180_o;
  wire n12182_o;
  wire [30:0] n12183_o;
  wire [31:0] n12184_o;
  wire n12186_o;
  wire n12187_o;
  wire n12188_o;
  wire n12190_o;
  wire [30:0] n12191_o;
  wire [31:0] n12192_o;
  wire n12194_o;
  wire n12195_o;
  wire n12197_o;
  wire n12201_o;
  wire n12202_o;
  wire n12203_o;
  wire n12206_o;
  wire [2:0] n12208_o;
  wire [2:0] n12209_o;
  wire [2:0] n12210_o;
  wire [5:0] n12211_o;
  wire [8:0] n12212_o;
  wire [2:0] n12213_o;
  wire [5:0] n12214_o;
  wire [5:0] n12215_o;
  wire [11:0] n12216_o;
  assign bus_addr_out = gen_src_addr_in;
  assign bus_addr_mode_out = gen_src_addr_mode_in;
  assign bus_cs_out = n12127_o;
  assign bus_read_out = n12129_o;
  assign bus_read_vm_out = gen_vm_in;
  assign bus_read_fork_out = gen_fork_in;
  assign bus_read_data_flow_out = gen_data_flow_in;
  assign bus_read_stream_out = gen_src_stream_in;
  assign bus_read_stream_id_out = gen_stream_id_in;
  assign bus_read_vector_out = gen_src_vector_in;
  assign bus_read_scatter_out = gen_src_scatter_in;
  assign bus_read_start_out = gen_src_start_in;
  assign bus_read_end_out = gen_src_end_in;
  assign bus_burstlen_out = gen_src_burstlen_in;
  assign bus_id_out = gen_bus_id_source_in;
  assign bus_data_type_out = gen_data_type_source_in;
  assign bus_data_model_out = gen_data_model_source_in;
  assign gen_waitreq_out = n12124_o;
  assign wr_req_out = n12208_o;
  assign wr_req_pending_p0_out = n12209_o;
  assign wr_req_pending_p1_out = n12210_o;
  assign wr_data_flow_out = n12211_o;
  assign wr_vector_out = n12212_o;
  assign wr_stream_out = n12213_o;
  assign wr_stream_id_out = n12214_o;
  assign wr_scatter_out = n12215_o;
  assign wr_end_out = n12216_o;
  assign wr_addr_out = wr_addr;
  assign wr_fork_out = wr_fork;
  assign wr_addr_mode_out = wr_addr_mode;
  assign wr_src_vm_out = wr_src_vm;
  assign wr_datavalid_out = n12132_o;
  assign wr_data_out = gen_src_data_in;
  assign wr_readdatavalid_out = bus_readdatavalid_in;
  assign wr_readdatavalid_vm_out = bus_readdatavalid_vm_in;
  assign wr_readdata_out = bus_readdata;
  assign wr_burstlen_out = wr_burstlen;
  assign wr_bus_id_out = dp_bus_id;
  assign wr_thread_out = dp_thread;
  assign wr_data_type_out = dp_data_type;
  assign wr_data_model_out = dp_data_model;
  assign wr_mcast_out = dp_mcast;
  /* ../../HW/src/dp/dp_source.vhd:135:8  */
  assign doit = gen_valid; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:136:8  */
  assign wr_req = n12206_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:137:8  */
  assign wr_addr = gen_dst_addr_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:138:8  */
  assign wr_fork = gen_fork_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:139:8  */
  assign wr_addr_mode = gen_dst_addr_mode_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:140:8  */
  assign wr_src_vm = gen_vm_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:141:8  */
  assign dp_bus_id = gen_bus_id_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:142:8  */
  assign dp_data_type = gen_data_type_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:143:8  */
  assign dp_data_model = gen_data_model_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:144:8  */
  assign dp_thread = gen_thread_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:145:8  */
  assign dp_mcast = gen_mcast_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:146:8  */
  assign wr_burstlen = gen_dst_burstlen_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:155:8  */
  assign gen_valid = n12078_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:156:8  */
  assign bus_readdata = n12079_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:160:32  */
  assign n12077_o = ~gen_busy_dest_in;
  /* ../../HW/src/dp/dp_source.vhd:160:27  */
  assign n12078_o = gen_valid_in & n12077_o;
  /* ../../HW/src/dp/dp_source.vhd:162:33  */
  assign n12079_o = bus_readdatavalid_in ? bus_readdata_in : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/dp/dp_source.vhd:164:1  */
  delay_8 delay_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_req),
    .enable_in(n12082_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:166:1  */
  delayi_2_8 delay_i3 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_bus_id),
    .enable_in(n12086_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:168:1  */
  delayi_2_8 delay_i4 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_data_type),
    .enable_in(n12090_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:170:1  */
  delayi_1_8 delay_i5 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_thread),
    .enable_in(n12094_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:172:1  */
  delayi_5_8 delay_i6 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_burstlen),
    .enable_in(n12098_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:174:1  */
  delayv_6_8 delay_i7 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_mcast),
    .enable_in(n12102_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:176:1  */
  delay_8 delay_i8 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(gen_src_eof_in),
    .enable_in(n12106_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:178:1  */
  delayv_64_8 delay_i9 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(gen_src_data_in),
    .enable_in(n12110_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:182:1  */
  delayv_64_4 gen_delay_i10 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(bus_readdata),
    .enable_in(n12114_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:190:39  */
  assign n12118_o = bus_wait_request_in & doit;
  /* ../../HW/src/dp/dp_source.vhd:190:85  */
  assign n12119_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:190:67  */
  assign n12120_o = n12119_o & n12118_o;
  /* ../../HW/src/dp/dp_source.vhd:190:104  */
  assign n12121_o = ~gen_valid;
  /* ../../HW/src/dp/dp_source.vhd:190:109  */
  assign n12122_o = gen_valid_in & n12121_o;
  /* ../../HW/src/dp/dp_source.vhd:190:91  */
  assign n12123_o = n12120_o | n12122_o;
  /* ../../HW/src/dp/dp_source.vhd:190:24  */
  assign n12124_o = n12123_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:202:30  */
  assign n12126_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:202:25  */
  assign n12127_o = gen_valid & n12126_o;
  /* ../../HW/src/dp/dp_source.vhd:203:32  */
  assign n12128_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:203:27  */
  assign n12129_o = gen_valid & n12128_o;
  /* ../../HW/src/dp/dp_source.vhd:234:21  */
  assign n12132_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n12135_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12136_o = {1'b0, n12135_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12138_o = 32'b00000000000000000000000000000000 == n12136_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12140_o = n12138_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12141_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12142_o = {1'b0, n12141_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12144_o = 32'b00000000000000000000000000000000 == n12142_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12145_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12146_o = gen_valid_in & n12145_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12148_o = n12144_o ? n12146_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12149_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12150_o = {1'b0, n12149_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12152_o = 32'b00000000000000000000000000000000 == n12150_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12153_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12155_o = n12152_o ? n12153_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n12156_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12157_o = {1'b0, n12156_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12159_o = 32'b00000000000000000000000000000001 == n12157_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12161_o = n12159_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12162_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12163_o = {1'b0, n12162_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12165_o = 32'b00000000000000000000000000000001 == n12163_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12166_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12167_o = gen_valid_in & n12166_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12169_o = n12165_o ? n12167_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12170_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12171_o = {1'b0, n12170_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12173_o = 32'b00000000000000000000000000000001 == n12171_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12174_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12176_o = n12173_o ? n12174_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n12177_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12178_o = {1'b0, n12177_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n12180_o = 32'b00000000000000000000000000000010 == n12178_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12182_o = n12180_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12183_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12184_o = {1'b0, n12183_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12186_o = 32'b00000000000000000000000000000010 == n12184_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12187_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12188_o = gen_valid_in & n12187_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12190_o = n12186_o ? n12188_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12191_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12192_o = {1'b0, n12191_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12194_o = 32'b00000000000000000000000000000010 == n12192_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12195_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12197_o = n12194_o ? n12195_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:278:41  */
  assign n12201_o = ~bus_wait_request_in;
  /* ../../HW/src/dp/dp_source.vhd:278:46  */
  assign n12202_o = n12201_o | gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:278:17  */
  assign n12203_o = n12202_o & doit;
  /* ../../HW/src/dp/dp_source.vhd:278:5  */
  assign n12206_o = n12203_o ? 1'b1 : 1'b0;
  assign n12208_o = {n12182_o, n12161_o, n12140_o};
  assign n12209_o = {n12190_o, n12169_o, n12148_o};
  assign n12210_o = {n12197_o, n12176_o, n12155_o};
  assign n12211_o = {gen_data_flow_in, gen_data_flow_in, gen_data_flow_in};
  assign n12212_o = {gen_dst_vector_in, gen_dst_vector_in, gen_dst_vector_in};
  assign n12213_o = {gen_dest_stream_in, gen_dest_stream_in, gen_dest_stream_in};
  assign n12214_o = {gen_stream_id_in, gen_stream_id_in, gen_stream_id_in};
  assign n12215_o = {gen_dst_scatter_in, gen_dst_scatter_in, gen_dst_scatter_in};
  assign n12216_o = {gen_dst_end_in, gen_dst_end_in, gen_dst_end_in};
endmodule

module dp_source_0_3_8_32_1_0
  (input  clock_in,
   input  reset_in,
   input  bus_readdatavalid_in,
   input  bus_readdatavalid_vm_in,
   input  [63:0] bus_readdata_in,
   input  bus_wait_request_in,
   input  gen_valid_in,
   input  gen_vm_in,
   input  gen_fork_in,
   input  [1:0] gen_data_flow_in,
   input  gen_src_stream_in,
   input  gen_dest_stream_in,
   input  [1:0] gen_stream_id_in,
   input  [2:0] gen_src_vector_in,
   input  [2:0] gen_dst_vector_in,
   input  [1:0] gen_src_scatter_in,
   input  [1:0] gen_dst_scatter_in,
   input  [3:0] gen_src_start_in,
   input  [3:0] gen_src_end_in,
   input  [3:0] gen_dst_end_in,
   input  gen_src_eof_in,
   input  [31:0] gen_src_addr_in,
   input  gen_src_addr_mode_in,
   input  [31:0] gen_dst_addr_in,
   input  gen_dst_addr_mode_in,
   input  [1:0] gen_bus_id_source_in,
   input  [1:0] gen_data_type_source_in,
   input  [1:0] gen_data_model_source_in,
   input  [1:0] gen_bus_id_dest_in,
   input  gen_busy_dest_in,
   input  [1:0] gen_data_type_dest_in,
   input  [1:0] gen_data_model_dest_in,
   input  [4:0] gen_src_burstlen_in,
   input  [4:0] gen_dst_burstlen_in,
   input  gen_thread_in,
   input  [5:0] gen_mcast_in,
   input  [63:0] gen_src_data_in,
   input  [2:0] wr_full_in,
   output [31:0] bus_addr_out,
   output bus_addr_mode_out,
   output bus_cs_out,
   output bus_read_out,
   output bus_read_vm_out,
   output bus_read_fork_out,
   output [1:0] bus_read_data_flow_out,
   output bus_read_stream_out,
   output [1:0] bus_read_stream_id_out,
   output [2:0] bus_read_vector_out,
   output [1:0] bus_read_scatter_out,
   output [3:0] bus_read_start_out,
   output [3:0] bus_read_end_out,
   output [4:0] bus_burstlen_out,
   output [1:0] bus_id_out,
   output [1:0] bus_data_type_out,
   output [1:0] bus_data_model_out,
   output gen_waitreq_out,
   output [2:0] wr_req_out,
   output [2:0] wr_req_pending_p0_out,
   output [2:0] wr_req_pending_p1_out,
   output [5:0] wr_data_flow_out,
   output [8:0] wr_vector_out,
   output [2:0] wr_stream_out,
   output [5:0] wr_stream_id_out,
   output [5:0] wr_scatter_out,
   output [11:0] wr_end_out,
   output [31:0] wr_addr_out,
   output wr_fork_out,
   output wr_addr_mode_out,
   output wr_src_vm_out,
   output wr_datavalid_out,
   output [63:0] wr_data_out,
   output wr_readdatavalid_out,
   output wr_readdatavalid_vm_out,
   output [63:0] wr_readdata_out,
   output [4:0] wr_burstlen_out,
   output [1:0] wr_bus_id_out,
   output wr_thread_out,
   output [1:0] wr_data_type_out,
   output [1:0] wr_data_model_out,
   output [5:0] wr_mcast_out);
  wire doit;
  wire wr_req;
  wire [31:0] wr_addr;
  wire wr_fork;
  wire wr_addr_mode;
  wire wr_src_vm;
  wire [1:0] dp_bus_id;
  wire [1:0] dp_data_type;
  wire [1:0] dp_data_model;
  wire dp_thread;
  wire [5:0] dp_mcast;
  wire [4:0] wr_burstlen;
  wire gen_valid;
  wire [63:0] bus_readdata;
  wire n11899_o;
  wire n11900_o;
  wire [63:0] n11901_o;
  localparam n11904_o = 1'b1;
  wire delay_i1_out_out;
  localparam n11908_o = 1'b1;
  wire [1:0] delay_i3_out_out;
  localparam n11912_o = 1'b1;
  wire [1:0] delay_i4_out_out;
  localparam n11916_o = 1'b1;
  wire delay_i5_out_out;
  localparam n11920_o = 1'b1;
  wire [4:0] delay_i6_out_out;
  localparam n11924_o = 1'b1;
  wire [5:0] delay_i7_out_out;
  localparam n11928_o = 1'b1;
  wire delay_i8_out_out;
  localparam n11932_o = 1'b1;
  wire [63:0] delay_i9_out_out;
  wire n11936_o;
  wire n11937_o;
  wire n11938_o;
  wire n11939_o;
  wire n11940_o;
  wire n11941_o;
  wire n11942_o;
  wire n11944_o;
  wire n11945_o;
  wire n11946_o;
  wire n11947_o;
  wire n11950_o;
  wire [30:0] n11953_o;
  wire [31:0] n11954_o;
  wire n11956_o;
  wire n11958_o;
  wire [30:0] n11959_o;
  wire [31:0] n11960_o;
  wire n11962_o;
  wire n11963_o;
  wire n11964_o;
  wire n11966_o;
  wire [30:0] n11967_o;
  wire [31:0] n11968_o;
  wire n11970_o;
  wire n11971_o;
  wire n11973_o;
  wire [30:0] n11974_o;
  wire [31:0] n11975_o;
  wire n11977_o;
  wire n11979_o;
  wire [30:0] n11980_o;
  wire [31:0] n11981_o;
  wire n11983_o;
  wire n11984_o;
  wire n11985_o;
  wire n11987_o;
  wire [30:0] n11988_o;
  wire [31:0] n11989_o;
  wire n11991_o;
  wire n11992_o;
  wire n11994_o;
  wire [30:0] n11995_o;
  wire [31:0] n11996_o;
  wire n11998_o;
  wire n12000_o;
  wire [30:0] n12001_o;
  wire [31:0] n12002_o;
  wire n12004_o;
  wire n12005_o;
  wire n12006_o;
  wire n12008_o;
  wire [30:0] n12009_o;
  wire [31:0] n12010_o;
  wire n12012_o;
  wire n12013_o;
  wire n12015_o;
  wire n12019_o;
  wire n12020_o;
  wire n12021_o;
  wire n12024_o;
  wire [2:0] n12026_o;
  wire [2:0] n12027_o;
  wire [2:0] n12028_o;
  wire [5:0] n12029_o;
  wire [8:0] n12030_o;
  wire [2:0] n12031_o;
  wire [5:0] n12032_o;
  wire [5:0] n12033_o;
  wire [11:0] n12034_o;
  assign bus_addr_out = gen_src_addr_in;
  assign bus_addr_mode_out = gen_src_addr_mode_in;
  assign bus_cs_out = n11945_o;
  assign bus_read_out = n11947_o;
  assign bus_read_vm_out = gen_vm_in;
  assign bus_read_fork_out = gen_fork_in;
  assign bus_read_data_flow_out = gen_data_flow_in;
  assign bus_read_stream_out = gen_src_stream_in;
  assign bus_read_stream_id_out = gen_stream_id_in;
  assign bus_read_vector_out = gen_src_vector_in;
  assign bus_read_scatter_out = gen_src_scatter_in;
  assign bus_read_start_out = gen_src_start_in;
  assign bus_read_end_out = gen_src_end_in;
  assign bus_burstlen_out = gen_src_burstlen_in;
  assign bus_id_out = gen_bus_id_source_in;
  assign bus_data_type_out = gen_data_type_source_in;
  assign bus_data_model_out = gen_data_model_source_in;
  assign gen_waitreq_out = n11942_o;
  assign wr_req_out = n12026_o;
  assign wr_req_pending_p0_out = n12027_o;
  assign wr_req_pending_p1_out = n12028_o;
  assign wr_data_flow_out = n12029_o;
  assign wr_vector_out = n12030_o;
  assign wr_stream_out = n12031_o;
  assign wr_stream_id_out = n12032_o;
  assign wr_scatter_out = n12033_o;
  assign wr_end_out = n12034_o;
  assign wr_addr_out = wr_addr;
  assign wr_fork_out = wr_fork;
  assign wr_addr_mode_out = wr_addr_mode;
  assign wr_src_vm_out = wr_src_vm;
  assign wr_datavalid_out = n11950_o;
  assign wr_data_out = gen_src_data_in;
  assign wr_readdatavalid_out = bus_readdatavalid_in;
  assign wr_readdatavalid_vm_out = bus_readdatavalid_vm_in;
  assign wr_readdata_out = bus_readdata;
  assign wr_burstlen_out = wr_burstlen;
  assign wr_bus_id_out = dp_bus_id;
  assign wr_thread_out = dp_thread;
  assign wr_data_type_out = dp_data_type;
  assign wr_data_model_out = dp_data_model;
  assign wr_mcast_out = dp_mcast;
  /* ../../HW/src/dp/dp_source.vhd:135:8  */
  assign doit = gen_valid; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:136:8  */
  assign wr_req = n12024_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:137:8  */
  assign wr_addr = gen_dst_addr_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:138:8  */
  assign wr_fork = gen_fork_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:139:8  */
  assign wr_addr_mode = gen_dst_addr_mode_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:140:8  */
  assign wr_src_vm = gen_vm_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:141:8  */
  assign dp_bus_id = gen_bus_id_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:142:8  */
  assign dp_data_type = gen_data_type_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:143:8  */
  assign dp_data_model = gen_data_model_dest_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:144:8  */
  assign dp_thread = gen_thread_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:145:8  */
  assign dp_mcast = gen_mcast_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:146:8  */
  assign wr_burstlen = gen_dst_burstlen_in; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:155:8  */
  assign gen_valid = n11900_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:156:8  */
  assign bus_readdata = n11901_o; // (signal)
  /* ../../HW/src/dp/dp_source.vhd:160:32  */
  assign n11899_o = ~gen_busy_dest_in;
  /* ../../HW/src/dp/dp_source.vhd:160:27  */
  assign n11900_o = gen_valid_in & n11899_o;
  /* ../../HW/src/dp/dp_source.vhd:162:33  */
  assign n11901_o = bus_readdatavalid_in ? bus_readdata_in : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/dp/dp_source.vhd:164:1  */
  delay_8 delay_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_req),
    .enable_in(n11904_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:166:1  */
  delayi_2_8 delay_i3 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_bus_id),
    .enable_in(n11908_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:168:1  */
  delayi_2_8 delay_i4 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_data_type),
    .enable_in(n11912_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:170:1  */
  delayi_1_8 delay_i5 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_thread),
    .enable_in(n11916_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:172:1  */
  delayi_5_8 delay_i6 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(wr_burstlen),
    .enable_in(n11920_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:174:1  */
  delayv_6_8 delay_i7 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(dp_mcast),
    .enable_in(n11924_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:176:1  */
  delay_8 delay_i8 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(gen_src_eof_in),
    .enable_in(n11928_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:178:1  */
  delayv_64_8 delay_i9 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(gen_src_data_in),
    .enable_in(n11932_o),
    .out_out());
  /* ../../HW/src/dp/dp_source.vhd:190:39  */
  assign n11936_o = bus_wait_request_in & doit;
  /* ../../HW/src/dp/dp_source.vhd:190:85  */
  assign n11937_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:190:67  */
  assign n11938_o = n11937_o & n11936_o;
  /* ../../HW/src/dp/dp_source.vhd:190:104  */
  assign n11939_o = ~gen_valid;
  /* ../../HW/src/dp/dp_source.vhd:190:109  */
  assign n11940_o = gen_valid_in & n11939_o;
  /* ../../HW/src/dp/dp_source.vhd:190:91  */
  assign n11941_o = n11938_o | n11940_o;
  /* ../../HW/src/dp/dp_source.vhd:190:24  */
  assign n11942_o = n11941_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:202:30  */
  assign n11944_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:202:25  */
  assign n11945_o = gen_valid & n11944_o;
  /* ../../HW/src/dp/dp_source.vhd:203:32  */
  assign n11946_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:203:27  */
  assign n11947_o = gen_valid & n11946_o;
  /* ../../HW/src/dp/dp_source.vhd:234:21  */
  assign n11950_o = ~gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n11953_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n11954_o = {1'b0, n11953_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n11956_o = 32'b00000000000000000000000000000000 == n11954_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n11958_o = n11956_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n11959_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n11960_o = {1'b0, n11959_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n11962_o = 32'b00000000000000000000000000000000 == n11960_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n11963_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n11964_o = gen_valid_in & n11963_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n11966_o = n11962_o ? n11964_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n11967_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n11968_o = {1'b0, n11967_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n11970_o = 32'b00000000000000000000000000000000 == n11968_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n11971_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n11973_o = n11970_o ? n11971_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n11974_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n11975_o = {1'b0, n11974_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n11977_o = 32'b00000000000000000000000000000001 == n11975_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n11979_o = n11977_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n11980_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n11981_o = {1'b0, n11980_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n11983_o = 32'b00000000000000000000000000000001 == n11981_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n11984_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n11985_o = gen_valid_in & n11984_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n11987_o = n11983_o ? n11985_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n11988_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n11989_o = {1'b0, n11988_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n11991_o = 32'b00000000000000000000000000000001 == n11989_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n11992_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n11994_o = n11991_o ? n11992_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:250:10  */
  assign n11995_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n11996_o = {1'b0, n11995_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:250:9  */
  assign n11998_o = 32'b00000000000000000000000000000010 == n11996_o;
  /* ../../HW/src/dp/dp_source.vhd:250:5  */
  assign n12000_o = n11998_o ? wr_req : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:255:10  */
  assign n12001_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12002_o = {1'b0, n12001_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:255:9  */
  assign n12004_o = 32'b00000000000000000000000000000010 == n12002_o;
  /* ../../HW/src/dp/dp_source.vhd:256:55  */
  assign n12005_o = ~gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:256:50  */
  assign n12006_o = gen_valid_in & n12005_o;
  /* ../../HW/src/dp/dp_source.vhd:255:5  */
  assign n12008_o = n12004_o ? n12006_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:260:10  */
  assign n12009_o = {29'b0, dp_bus_id};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12010_o = {1'b0, n12009_o};  //  uext
  /* ../../HW/src/dp/dp_source.vhd:260:9  */
  assign n12012_o = 32'b00000000000000000000000000000010 == n12010_o;
  /* ../../HW/src/dp/dp_source.vhd:261:50  */
  assign n12013_o = gen_valid_in & gen_vm_in;
  /* ../../HW/src/dp/dp_source.vhd:260:5  */
  assign n12015_o = n12012_o ? n12013_o : 1'b0;
  /* ../../HW/src/dp/dp_source.vhd:278:41  */
  assign n12019_o = ~bus_wait_request_in;
  /* ../../HW/src/dp/dp_source.vhd:278:46  */
  assign n12020_o = n12019_o | gen_src_eof_in;
  /* ../../HW/src/dp/dp_source.vhd:278:17  */
  assign n12021_o = n12020_o & doit;
  /* ../../HW/src/dp/dp_source.vhd:278:5  */
  assign n12024_o = n12021_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_gen_core.vhd:80:15  */
  assign n12026_o = {n12000_o, n11979_o, n11958_o};
  /* ../../HW/src/dp/dp_gen_core.vhd:79:15  */
  assign n12027_o = {n12008_o, n11987_o, n11966_o};
  /* ../../HW/src/dp/dp_gen_core.vhd:78:15  */
  assign n12028_o = {n12015_o, n11994_o, n11973_o};
  /* ../../HW/src/dp/dp_gen_core.vhd:77:15  */
  assign n12029_o = {gen_data_flow_in, gen_data_flow_in, gen_data_flow_in};
  /* ../../HW/src/dp/dp_gen_core.vhd:76:15  */
  assign n12030_o = {gen_dst_vector_in, gen_dst_vector_in, gen_dst_vector_in};
  /* ../../HW/src/dp/dp_gen_core.vhd:75:15  */
  assign n12031_o = {gen_dest_stream_in, gen_dest_stream_in, gen_dest_stream_in};
  /* ../../HW/src/dp/dp_gen_core.vhd:74:15  */
  assign n12032_o = {gen_stream_id_in, gen_stream_id_in, gen_stream_id_in};
  /* ../../HW/src/dp/dp_gen_core.vhd:73:15  */
  assign n12033_o = {gen_dst_scatter_in, gen_dst_scatter_in, gen_dst_scatter_in};
  /* ../../HW/src/dp/dp_gen_core.vhd:72:15  */
  assign n12034_o = {gen_dst_end_in, gen_dst_end_in, gen_dst_end_in};
endmodule

module dp_gen_core
  (input  clock_in,
   input  reset_in,
   input  [1:0] instruction_valid_in,
   input  [2:0] instruction_in_opcode,
   input  [3:0] instruction_in_condition,
   input  instruction_in_vm,
   input  [775:0] instruction_in_source,
   input  [1:0] instruction_in_source_bus_id,
   input  [1:0] instruction_in_source_data_type,
   input  [775:0] instruction_in_dest,
   input  [1:0] instruction_in_dest_bus_id,
   input  [1:0] instruction_in_dest_data_type,
   input  [5:0] instruction_in_mcast,
   input  [23:0] instruction_in_count,
   input  [15:0] instruction_in_data,
   input  instruction_in_repeat,
   input  instruction_in_source_addr_mode,
   input  instruction_in_dest_addr_mode,
   input  instruction_in_stream_process,
   input  [1:0] instruction_in_stream_process_id,
   input  [2:0] pre_instruction_in_opcode,
   input  [3:0] pre_instruction_in_condition,
   input  pre_instruction_in_vm,
   input  [775:0] pre_instruction_in_source,
   input  [1:0] pre_instruction_in_source_bus_id,
   input  [1:0] pre_instruction_in_source_data_type,
   input  [775:0] pre_instruction_in_dest,
   input  [1:0] pre_instruction_in_dest_bus_id,
   input  [1:0] pre_instruction_in_dest_data_type,
   input  [5:0] pre_instruction_in_mcast,
   input  [23:0] pre_instruction_in_count,
   input  [15:0] pre_instruction_in_data,
   input  pre_instruction_in_repeat,
   input  pre_instruction_in_source_addr_mode,
   input  pre_instruction_in_dest_addr_mode,
   input  pre_instruction_in_stream_process,
   input  [1:0] pre_instruction_in_stream_process_id,
   input  [14:0] wr_maxburstlen_in,
   input  [2:0] full_in,
   input  [2:0] waitreq_in,
   input  [71:0] bar_in,
   output [1:0] ready_out,
   output [31:0] log1_out,
   output log1_valid_out,
   output [31:0] log2_out,
   output log2_valid_out,
   output gen_pcore_src_valid_out,
   output gen_pcore_vm_out,
   output gen_pcore_fork_out,
   output [1:0] gen_pcore_data_flow_out,
   output gen_pcore_src_stream_out,
   output gen_pcore_dest_stream_out,
   output [1:0] gen_pcore_stream_id_out,
   output [2:0] gen_pcore_src_vector_out,
   output [2:0] gen_pcore_dst_vector_out,
   output [1:0] gen_pcore_src_scatter_out,
   output [1:0] gen_pcore_dst_scatter_out,
   output [3:0] gen_pcore_src_start_out,
   output [3:0] gen_pcore_src_end_out,
   output [3:0] gen_pcore_dst_end_out,
   output [31:0] gen_pcore_src_addr_out,
   output gen_pcore_src_addr_mode_out,
   output [31:0] gen_pcore_dst_addr_out,
   output gen_pcore_dst_addr_mode_out,
   output gen_pcore_src_eof_out,
   output [1:0] gen_pcore_bus_id_source_out,
   output [1:0] gen_pcore_data_type_source_out,
   output [1:0] gen_pcore_data_model_source_out,
   output [1:0] gen_pcore_bus_id_dest_out,
   output gen_pcore_busy_dest_out,
   output [1:0] gen_pcore_data_type_dest_out,
   output [1:0] gen_pcore_data_model_dest_out,
   output [4:0] gen_pcore_src_burstlen_out,
   output [4:0] gen_pcore_dst_burstlen_out,
   output gen_pcore_thread_out,
   output [5:0] gen_pcore_mcast_out,
   output [63:0] gen_pcore_data_out,
   output gen_sram_src_valid_out,
   output gen_sram_vm_out,
   output gen_sram_fork_out,
   output [1:0] gen_sram_data_flow_out,
   output gen_sram_src_stream_out,
   output gen_sram_dest_stream_out,
   output [1:0] gen_sram_stream_id_out,
   output [2:0] gen_sram_src_vector_out,
   output [2:0] gen_sram_dst_vector_out,
   output [1:0] gen_sram_src_scatter_out,
   output [1:0] gen_sram_dst_scatter_out,
   output [3:0] gen_sram_src_start_out,
   output [3:0] gen_sram_src_end_out,
   output [3:0] gen_sram_dst_end_out,
   output [31:0] gen_sram_src_addr_out,
   output gen_sram_src_addr_mode_out,
   output [31:0] gen_sram_dst_addr_out,
   output gen_sram_dst_addr_mode_out,
   output gen_sram_src_eof_out,
   output [1:0] gen_sram_bus_id_source_out,
   output [1:0] gen_sram_data_type_source_out,
   output [1:0] gen_sram_data_model_source_out,
   output [1:0] gen_sram_bus_id_dest_out,
   output gen_sram_busy_dest_out,
   output [1:0] gen_sram_data_type_dest_out,
   output [1:0] gen_sram_data_model_dest_out,
   output [4:0] gen_sram_src_burstlen_out,
   output [4:0] gen_sram_dst_burstlen_out,
   output gen_sram_thread_out,
   output [5:0] gen_sram_mcast_out,
   output [63:0] gen_sram_data_out,
   output gen_ddr_src_valid_out,
   output gen_ddr_vm_out,
   output gen_ddr_fork_out,
   output [1:0] gen_ddr_data_flow_out,
   output gen_ddr_src_stream_out,
   output gen_ddr_dest_stream_out,
   output [1:0] gen_ddr_stream_id_out,
   output [2:0] gen_ddr_src_vector_out,
   output [2:0] gen_ddr_dst_vector_out,
   output [1:0] gen_ddr_src_scatter_out,
   output [1:0] gen_ddr_dst_scatter_out,
   output [3:0] gen_ddr_src_start_out,
   output [3:0] gen_ddr_src_end_out,
   output [3:0] gen_ddr_dst_end_out,
   output [31:0] gen_ddr_src_addr_out,
   output gen_ddr_src_addr_mode_out,
   output [31:0] gen_ddr_dst_addr_out,
   output gen_ddr_dst_addr_mode_out,
   output gen_ddr_src_eof_out,
   output [1:0] gen_ddr_bus_id_source_out,
   output [1:0] gen_ddr_data_type_source_out,
   output [1:0] gen_ddr_data_model_source_out,
   output [1:0] gen_ddr_bus_id_dest_out,
   output gen_ddr_busy_dest_out,
   output [1:0] gen_ddr_data_type_dest_out,
   output [1:0] gen_ddr_data_model_dest_out,
   output [4:0] gen_ddr_src_burstlen_out,
   output [4:0] gen_ddr_dst_burstlen_out,
   output gen_ddr_thread_out,
   output [5:0] gen_ddr_mcast_out,
   output [63:0] gen_ddr_data_out);
  wire [1619:0] n11072_o;
  wire [1619:0] n11073_o;
  wire [2:0] gen_src_valid_1;
  wire gen_fork_1;
  wire gen_vm_1;
  wire [1:0] gen_data_flow_1;
  wire gen_src_stream_1;
  wire gen_dest_stream_1;
  wire [1:0] gen_stream_id_1;
  wire [2:0] gen_src_vector_1;
  wire [2:0] gen_dst_vector_1;
  wire [1:0] gen_src_scatter_1;
  wire [1:0] gen_dst_scatter_1;
  wire [3:0] gen_src_start_1;
  wire [3:0] gen_src_end_1;
  wire [3:0] gen_dst_end_1;
  wire [31:0] gen_src_addr_1;
  wire gen_src_addr_mode_1;
  wire [31:0] gen_dst_addr_1;
  wire gen_dst_addr_mode_1;
  wire gen_src_eof_1;
  wire [1:0] gen_bus_id_source_1;
  wire [1:0] gen_data_type_source_1;
  wire [1:0] gen_data_model_source_1;
  wire [1:0] gen_bus_id_dest_1;
  wire gen_busy_dest_1;
  wire [1:0] gen_data_type_dest_1;
  wire [1:0] gen_data_model_dest_1;
  wire [4:0] gen_src_burstlen_1;
  wire [4:0] gen_dst_burstlen_1;
  wire gen_thread_1;
  wire [5:0] gen_mcast_1;
  wire [63:0] gen_data_1;
  wire [2:0] gen_src_valid_2;
  wire gen_vm_2;
  wire gen_fork_2;
  wire [1:0] gen_data_flow_2;
  wire gen_src_stream_2;
  wire gen_dest_stream_2;
  wire [1:0] gen_stream_id_2;
  wire [2:0] gen_src_vector_2;
  wire [2:0] gen_dst_vector_2;
  wire [1:0] gen_src_scatter_2;
  wire [1:0] gen_dst_scatter_2;
  wire [3:0] gen_src_start_2;
  wire [3:0] gen_src_end_2;
  wire [3:0] gen_dst_end_2;
  wire [31:0] gen_src_addr_2;
  wire gen_src_addr_mode_2;
  wire [31:0] gen_dst_addr_2;
  wire gen_dst_addr_mode_2;
  wire gen_src_eof_2;
  wire [1:0] gen_bus_id_source_2;
  wire [1:0] gen_data_type_source_2;
  wire [1:0] gen_data_model_source_2;
  wire [1:0] gen_bus_id_dest_2;
  wire gen_busy_dest_2;
  wire [1:0] gen_data_type_dest_2;
  wire [1:0] gen_data_model_dest_2;
  wire [4:0] gen_src_burstlen_2;
  wire [4:0] gen_dst_burstlen_2;
  wire gen_thread_2;
  wire [5:0] gen_mcast_2;
  wire [63:0] gen_data_2;
  wire [1:0] ready;
  wire n11173_o;
  wire n11175_o;
  wire n11177_o;
  wire n11178_o;
  wire n11179_o;
  wire n11180_o;
  wire [1:0] n11181_o;
  wire n11182_o;
  wire n11183_o;
  wire [1:0] n11184_o;
  wire [2:0] n11185_o;
  wire [2:0] n11186_o;
  wire [1:0] n11187_o;
  wire [1:0] n11188_o;
  wire [3:0] n11189_o;
  wire [3:0] n11190_o;
  wire [3:0] n11191_o;
  wire [31:0] n11192_o;
  wire n11193_o;
  wire [31:0] n11194_o;
  wire n11195_o;
  wire n11196_o;
  wire [1:0] n11197_o;
  wire [1:0] n11198_o;
  wire [1:0] n11199_o;
  wire [1:0] n11200_o;
  wire n11201_o;
  wire [1:0] n11202_o;
  wire [1:0] n11203_o;
  wire [4:0] n11204_o;
  wire [4:0] n11205_o;
  wire n11206_o;
  wire [5:0] n11207_o;
  wire [63:0] n11208_o;
  wire n11213_o;
  wire n11214_o;
  wire n11215_o;
  wire n11216_o;
  wire n11217_o;
  wire n11218_o;
  wire [1:0] n11219_o;
  wire n11220_o;
  wire n11221_o;
  wire [1:0] n11222_o;
  wire [2:0] n11223_o;
  wire [2:0] n11224_o;
  wire [1:0] n11225_o;
  wire [1:0] n11226_o;
  wire [3:0] n11227_o;
  wire [3:0] n11228_o;
  wire [3:0] n11229_o;
  wire [31:0] n11230_o;
  wire n11231_o;
  wire [31:0] n11232_o;
  wire n11233_o;
  wire n11234_o;
  wire [1:0] n11235_o;
  wire [1:0] n11236_o;
  wire [1:0] n11237_o;
  wire [1:0] n11238_o;
  wire n11239_o;
  wire [1:0] n11240_o;
  wire [1:0] n11241_o;
  wire [4:0] n11242_o;
  wire [4:0] n11243_o;
  wire n11244_o;
  wire [5:0] n11245_o;
  wire [63:0] n11246_o;
  wire n11250_o;
  wire n11252_o;
  wire n11254_o;
  wire n11255_o;
  wire n11256_o;
  wire n11257_o;
  wire [1:0] n11258_o;
  wire n11259_o;
  wire n11260_o;
  wire [1:0] n11261_o;
  wire [2:0] n11262_o;
  wire [2:0] n11263_o;
  wire [1:0] n11264_o;
  wire [1:0] n11265_o;
  wire [3:0] n11266_o;
  wire [3:0] n11267_o;
  wire [3:0] n11268_o;
  wire [31:0] n11269_o;
  wire n11270_o;
  wire [31:0] n11271_o;
  wire n11272_o;
  wire n11273_o;
  wire [1:0] n11274_o;
  wire [1:0] n11275_o;
  wire [1:0] n11276_o;
  wire [1:0] n11277_o;
  wire n11278_o;
  wire [1:0] n11279_o;
  wire [1:0] n11280_o;
  wire [4:0] n11281_o;
  wire [4:0] n11282_o;
  wire n11283_o;
  wire [5:0] n11284_o;
  wire [63:0] n11285_o;
  wire dp_gen_primary_i_n11288;
  wire n11289_o;
  wire n11290_o;
  wire [775:0] n11291_o;
  wire [775:0] n11292_o;
  wire n11293_o;
  wire [1:0] n11294_o;
  wire n11295_o;
  wire [775:0] n11296_o;
  wire [775:0] n11297_o;
  wire [1:0] n11298_o;
  wire [1:0] n11299_o;
  wire n11300_o;
  wire n11301_o;
  wire [1:0] n11302_o;
  wire [1:0] n11303_o;
  wire [775:0] n11304_o;
  wire [1:0] n11305_o;
  wire [1:0] n11306_o;
  wire [1:0] n11307_o;
  wire [775:0] n11308_o;
  wire [1:0] n11309_o;
  wire [5:0] n11310_o;
  wire [23:0] n11311_o;
  localparam n11312_o = 1'b0;
  wire [15:0] n11313_o;
  wire n11314_o;
  wire [2:0] dp_gen_primary_i_n11315;
  wire dp_gen_primary_i_n11316;
  wire dp_gen_primary_i_n11317;
  wire [1:0] dp_gen_primary_i_n11318;
  wire dp_gen_primary_i_n11319;
  wire dp_gen_primary_i_n11320;
  wire [1:0] dp_gen_primary_i_n11321;
  wire [2:0] dp_gen_primary_i_n11322;
  wire [2:0] dp_gen_primary_i_n11323;
  wire [1:0] dp_gen_primary_i_n11324;
  wire [1:0] dp_gen_primary_i_n11325;
  wire [3:0] dp_gen_primary_i_n11326;
  wire [3:0] dp_gen_primary_i_n11327;
  wire [3:0] dp_gen_primary_i_n11328;
  wire [31:0] dp_gen_primary_i_n11329;
  wire dp_gen_primary_i_n11330;
  wire [31:0] dp_gen_primary_i_n11331;
  wire dp_gen_primary_i_n11332;
  wire dp_gen_primary_i_n11333;
  wire [1:0] dp_gen_primary_i_n11334;
  wire [1:0] dp_gen_primary_i_n11335;
  wire [1:0] dp_gen_primary_i_n11336;
  wire [1:0] dp_gen_primary_i_n11337;
  wire dp_gen_primary_i_n11338;
  wire [1:0] dp_gen_primary_i_n11339;
  wire [1:0] dp_gen_primary_i_n11340;
  wire [4:0] dp_gen_primary_i_n11341;
  wire [4:0] dp_gen_primary_i_n11342;
  wire dp_gen_primary_i_n11343;
  wire [5:0] dp_gen_primary_i_n11344;
  wire [63:0] dp_gen_primary_i_n11345;
  wire [31:0] dp_gen_primary_i_n11346;
  wire dp_gen_primary_i_n11347;
  wire dp_gen_primary_i_ready_out;
  wire [2:0] dp_gen_primary_i_gen_valid_out;
  wire dp_gen_primary_i_gen_vm_out;
  wire dp_gen_primary_i_gen_fork_out;
  wire [1:0] dp_gen_primary_i_gen_data_flow_out;
  wire dp_gen_primary_i_gen_src_stream_out;
  wire dp_gen_primary_i_gen_dest_stream_out;
  wire [1:0] dp_gen_primary_i_gen_stream_id_out;
  wire [2:0] dp_gen_primary_i_gen_src_vector_out;
  wire [2:0] dp_gen_primary_i_gen_dst_vector_out;
  wire [1:0] dp_gen_primary_i_gen_src_scatter_out;
  wire [1:0] dp_gen_primary_i_gen_dst_scatter_out;
  wire [3:0] dp_gen_primary_i_gen_src_start_out;
  wire [3:0] dp_gen_primary_i_gen_src_end_out;
  wire [3:0] dp_gen_primary_i_gen_dst_end_out;
  wire [31:0] dp_gen_primary_i_gen_addr_source_out;
  wire dp_gen_primary_i_gen_addr_source_mode_out;
  wire [31:0] dp_gen_primary_i_gen_addr_dest_out;
  wire dp_gen_primary_i_gen_addr_dest_mode_out;
  wire dp_gen_primary_i_gen_eof_out;
  wire [1:0] dp_gen_primary_i_gen_bus_id_source_out;
  wire [1:0] dp_gen_primary_i_gen_data_type_source_out;
  wire [1:0] dp_gen_primary_i_gen_data_model_source_out;
  wire [1:0] dp_gen_primary_i_gen_bus_id_dest_out;
  wire dp_gen_primary_i_gen_busy_dest_out;
  wire [1:0] dp_gen_primary_i_gen_data_type_dest_out;
  wire [1:0] dp_gen_primary_i_gen_data_model_dest_out;
  wire [4:0] dp_gen_primary_i_gen_burstlen_source_out;
  wire [4:0] dp_gen_primary_i_gen_burstlen_dest_out;
  wire dp_gen_primary_i_gen_thread_out;
  wire [5:0] dp_gen_primary_i_gen_mcast_out;
  wire [63:0] dp_gen_primary_i_gen_data_out;
  wire [31:0] dp_gen_primary_i_log_out;
  wire dp_gen_primary_i_log_valid_out;
  wire [23:0] n11349_o;
  wire [23:0] n11350_o;
  wire [24:0] n11351_o;
  wire [24:0] n11352_o;
  wire [23:0] n11353_o;
  wire [23:0] n11354_o;
  wire [24:0] n11355_o;
  wire [24:0] n11356_o;
  wire [23:0] n11357_o;
  wire [23:0] n11358_o;
  wire [24:0] n11359_o;
  wire [24:0] n11360_o;
  wire [23:0] n11361_o;
  wire [23:0] n11362_o;
  wire [24:0] n11363_o;
  wire [24:0] n11364_o;
  wire [23:0] n11365_o;
  wire [23:0] n11366_o;
  wire [24:0] n11367_o;
  wire [24:0] n11368_o;
  wire [24:0] n11369_o;
  wire [24:0] n11370_o;
  wire [24:0] n11371_o;
  wire [2:0] n11372_o;
  wire [24:0] n11373_o;
  wire [31:0] n11374_o;
  wire [23:0] n11375_o;
  wire [23:0] n11376_o;
  wire n11377_o;
  wire [1:0] n11378_o;
  wire n11379_o;
  wire [23:0] n11380_o;
  wire [5:0] n11381_o;
  wire [15:0] n11382_o;
  wire n11383_o;
  wire [1:0] n11384_o;
  wire [1:0] n11385_o;
  wire [23:0] n11386_o;
  wire [23:0] n11387_o;
  wire [23:0] n11388_o;
  wire [23:0] n11389_o;
  wire [24:0] n11390_o;
  wire [24:0] n11391_o;
  wire [23:0] n11392_o;
  wire [23:0] n11393_o;
  wire [24:0] n11394_o;
  wire [24:0] n11395_o;
  wire [23:0] n11396_o;
  wire [23:0] n11397_o;
  wire [24:0] n11398_o;
  wire [24:0] n11399_o;
  wire [23:0] n11400_o;
  wire [23:0] n11401_o;
  wire [24:0] n11402_o;
  wire [24:0] n11403_o;
  wire [23:0] n11404_o;
  wire [23:0] n11405_o;
  wire [24:0] n11406_o;
  wire [24:0] n11407_o;
  wire [24:0] n11408_o;
  wire [24:0] n11409_o;
  wire [24:0] n11410_o;
  wire [2:0] n11411_o;
  wire [24:0] n11412_o;
  wire [31:0] n11413_o;
  wire [23:0] n11414_o;
  wire [23:0] n11415_o;
  wire n11416_o;
  wire [1:0] n11417_o;
  wire n11418_o;
  wire [23:0] n11419_o;
  wire [5:0] n11420_o;
  wire [15:0] n11421_o;
  wire n11422_o;
  wire [1:0] n11423_o;
  wire [1:0] n11424_o;
  wire [23:0] n11425_o;
  wire [23:0] n11426_o;
  wire [23:0] n11427_o;
  wire [23:0] n11428_o;
  wire [24:0] n11429_o;
  wire [24:0] n11430_o;
  wire [23:0] n11431_o;
  wire [23:0] n11432_o;
  wire [24:0] n11433_o;
  wire [24:0] n11434_o;
  wire [23:0] n11435_o;
  wire [23:0] n11436_o;
  wire [24:0] n11437_o;
  wire [24:0] n11438_o;
  wire [23:0] n11439_o;
  wire [23:0] n11440_o;
  wire [24:0] n11441_o;
  wire [24:0] n11442_o;
  wire [23:0] n11443_o;
  wire [23:0] n11444_o;
  wire [24:0] n11445_o;
  wire [24:0] n11446_o;
  wire [24:0] n11447_o;
  wire [24:0] n11448_o;
  wire [24:0] n11449_o;
  wire [2:0] n11450_o;
  wire [24:0] n11451_o;
  wire [31:0] n11452_o;
  wire [23:0] n11453_o;
  wire [23:0] n11454_o;
  wire n11455_o;
  wire [1:0] n11456_o;
  wire n11457_o;
  wire [23:0] n11458_o;
  wire [5:0] n11459_o;
  wire [15:0] n11460_o;
  wire n11461_o;
  wire [1:0] n11462_o;
  wire [1:0] n11463_o;
  wire [23:0] n11464_o;
  wire [23:0] n11465_o;
  wire [23:0] n11466_o;
  wire [23:0] n11467_o;
  wire [24:0] n11468_o;
  wire [24:0] n11469_o;
  wire [23:0] n11470_o;
  wire [23:0] n11471_o;
  wire [24:0] n11472_o;
  wire [24:0] n11473_o;
  wire [23:0] n11474_o;
  wire [23:0] n11475_o;
  wire [24:0] n11476_o;
  wire [24:0] n11477_o;
  wire [23:0] n11478_o;
  wire [23:0] n11479_o;
  wire [24:0] n11480_o;
  wire [24:0] n11481_o;
  wire [23:0] n11482_o;
  wire [23:0] n11483_o;
  wire [24:0] n11484_o;
  wire [24:0] n11485_o;
  wire [24:0] n11486_o;
  wire [24:0] n11487_o;
  wire [24:0] n11488_o;
  wire [2:0] n11489_o;
  wire [24:0] n11490_o;
  wire [31:0] n11491_o;
  wire [23:0] n11492_o;
  wire [23:0] n11493_o;
  wire n11494_o;
  wire [1:0] n11495_o;
  wire n11496_o;
  wire [23:0] n11497_o;
  wire [5:0] n11498_o;
  wire [15:0] n11499_o;
  wire n11500_o;
  wire [1:0] n11501_o;
  wire [1:0] n11502_o;
  wire [23:0] n11503_o;
  wire [23:0] n11504_o;
  wire dp_gen_secondary_i_n11572;
  wire n11573_o;
  wire n11574_o;
  wire [775:0] n11575_o;
  wire [775:0] n11576_o;
  wire n11577_o;
  wire [1:0] n11578_o;
  wire n11579_o;
  wire [775:0] n11580_o;
  wire [775:0] n11581_o;
  wire [1:0] n11582_o;
  wire [1:0] n11583_o;
  wire n11584_o;
  wire n11585_o;
  wire [1:0] n11586_o;
  wire [1:0] n11587_o;
  wire [775:0] n11588_o;
  wire [1:0] n11589_o;
  wire [1:0] n11590_o;
  wire [1:0] n11591_o;
  wire [775:0] n11592_o;
  wire [1:0] n11593_o;
  wire [5:0] n11594_o;
  wire [23:0] n11595_o;
  localparam n11596_o = 1'b0;
  wire [15:0] n11597_o;
  wire n11598_o;
  wire [2:0] dp_gen_secondary_i_n11599;
  wire dp_gen_secondary_i_n11600;
  wire dp_gen_secondary_i_n11601;
  wire [1:0] dp_gen_secondary_i_n11602;
  wire dp_gen_secondary_i_n11603;
  wire dp_gen_secondary_i_n11604;
  wire [1:0] dp_gen_secondary_i_n11605;
  wire [2:0] dp_gen_secondary_i_n11606;
  wire [2:0] dp_gen_secondary_i_n11607;
  wire [1:0] dp_gen_secondary_i_n11608;
  wire [1:0] dp_gen_secondary_i_n11609;
  wire [3:0] dp_gen_secondary_i_n11610;
  wire [3:0] dp_gen_secondary_i_n11611;
  wire [3:0] dp_gen_secondary_i_n11612;
  wire [31:0] dp_gen_secondary_i_n11613;
  wire dp_gen_secondary_i_n11614;
  wire [31:0] dp_gen_secondary_i_n11615;
  wire dp_gen_secondary_i_n11616;
  wire dp_gen_secondary_i_n11617;
  wire [1:0] dp_gen_secondary_i_n11618;
  wire [1:0] dp_gen_secondary_i_n11619;
  wire [1:0] dp_gen_secondary_i_n11620;
  wire [1:0] dp_gen_secondary_i_n11621;
  wire dp_gen_secondary_i_n11622;
  wire [1:0] dp_gen_secondary_i_n11623;
  wire [1:0] dp_gen_secondary_i_n11624;
  wire [4:0] dp_gen_secondary_i_n11625;
  wire [4:0] dp_gen_secondary_i_n11626;
  wire dp_gen_secondary_i_n11627;
  wire [5:0] dp_gen_secondary_i_n11628;
  wire [63:0] dp_gen_secondary_i_n11629;
  wire [31:0] dp_gen_secondary_i_n11630;
  wire dp_gen_secondary_i_n11631;
  wire dp_gen_secondary_i_ready_out;
  wire [2:0] dp_gen_secondary_i_gen_valid_out;
  wire dp_gen_secondary_i_gen_vm_out;
  wire dp_gen_secondary_i_gen_fork_out;
  wire [1:0] dp_gen_secondary_i_gen_data_flow_out;
  wire dp_gen_secondary_i_gen_src_stream_out;
  wire dp_gen_secondary_i_gen_dest_stream_out;
  wire [1:0] dp_gen_secondary_i_gen_stream_id_out;
  wire [2:0] dp_gen_secondary_i_gen_src_vector_out;
  wire [2:0] dp_gen_secondary_i_gen_dst_vector_out;
  wire [1:0] dp_gen_secondary_i_gen_src_scatter_out;
  wire [1:0] dp_gen_secondary_i_gen_dst_scatter_out;
  wire [3:0] dp_gen_secondary_i_gen_src_start_out;
  wire [3:0] dp_gen_secondary_i_gen_src_end_out;
  wire [3:0] dp_gen_secondary_i_gen_dst_end_out;
  wire [31:0] dp_gen_secondary_i_gen_addr_source_out;
  wire dp_gen_secondary_i_gen_addr_source_mode_out;
  wire [31:0] dp_gen_secondary_i_gen_addr_dest_out;
  wire dp_gen_secondary_i_gen_addr_dest_mode_out;
  wire dp_gen_secondary_i_gen_eof_out;
  wire [1:0] dp_gen_secondary_i_gen_bus_id_source_out;
  wire [1:0] dp_gen_secondary_i_gen_data_type_source_out;
  wire [1:0] dp_gen_secondary_i_gen_data_model_source_out;
  wire [1:0] dp_gen_secondary_i_gen_bus_id_dest_out;
  wire dp_gen_secondary_i_gen_busy_dest_out;
  wire [1:0] dp_gen_secondary_i_gen_data_type_dest_out;
  wire [1:0] dp_gen_secondary_i_gen_data_model_dest_out;
  wire [4:0] dp_gen_secondary_i_gen_burstlen_source_out;
  wire [4:0] dp_gen_secondary_i_gen_burstlen_dest_out;
  wire dp_gen_secondary_i_gen_thread_out;
  wire [5:0] dp_gen_secondary_i_gen_mcast_out;
  wire [63:0] dp_gen_secondary_i_gen_data_out;
  wire [31:0] dp_gen_secondary_i_log_out;
  wire dp_gen_secondary_i_log_valid_out;
  wire [23:0] n11633_o;
  wire [23:0] n11634_o;
  wire [24:0] n11635_o;
  wire [24:0] n11636_o;
  wire [23:0] n11637_o;
  wire [23:0] n11638_o;
  wire [24:0] n11639_o;
  wire [24:0] n11640_o;
  wire [23:0] n11641_o;
  wire [23:0] n11642_o;
  wire [24:0] n11643_o;
  wire [24:0] n11644_o;
  wire [23:0] n11645_o;
  wire [23:0] n11646_o;
  wire [24:0] n11647_o;
  wire [24:0] n11648_o;
  wire [23:0] n11649_o;
  wire [23:0] n11650_o;
  wire [24:0] n11651_o;
  wire [24:0] n11652_o;
  wire [24:0] n11653_o;
  wire [24:0] n11654_o;
  wire [24:0] n11655_o;
  wire [2:0] n11656_o;
  wire [24:0] n11657_o;
  wire [31:0] n11658_o;
  wire [23:0] n11659_o;
  wire [23:0] n11660_o;
  wire n11661_o;
  wire [1:0] n11662_o;
  wire n11663_o;
  wire [23:0] n11664_o;
  wire [5:0] n11665_o;
  wire [15:0] n11666_o;
  wire n11667_o;
  wire [1:0] n11668_o;
  wire [1:0] n11669_o;
  wire [23:0] n11670_o;
  wire [23:0] n11671_o;
  wire [23:0] n11672_o;
  wire [23:0] n11673_o;
  wire [24:0] n11674_o;
  wire [24:0] n11675_o;
  wire [23:0] n11676_o;
  wire [23:0] n11677_o;
  wire [24:0] n11678_o;
  wire [24:0] n11679_o;
  wire [23:0] n11680_o;
  wire [23:0] n11681_o;
  wire [24:0] n11682_o;
  wire [24:0] n11683_o;
  wire [23:0] n11684_o;
  wire [23:0] n11685_o;
  wire [24:0] n11686_o;
  wire [24:0] n11687_o;
  wire [23:0] n11688_o;
  wire [23:0] n11689_o;
  wire [24:0] n11690_o;
  wire [24:0] n11691_o;
  wire [24:0] n11692_o;
  wire [24:0] n11693_o;
  wire [24:0] n11694_o;
  wire [2:0] n11695_o;
  wire [24:0] n11696_o;
  wire [31:0] n11697_o;
  wire [23:0] n11698_o;
  wire [23:0] n11699_o;
  wire n11700_o;
  wire [1:0] n11701_o;
  wire n11702_o;
  wire [23:0] n11703_o;
  wire [5:0] n11704_o;
  wire [15:0] n11705_o;
  wire n11706_o;
  wire [1:0] n11707_o;
  wire [1:0] n11708_o;
  wire [23:0] n11709_o;
  wire [23:0] n11710_o;
  wire [23:0] n11711_o;
  wire [23:0] n11712_o;
  wire [24:0] n11713_o;
  wire [24:0] n11714_o;
  wire [23:0] n11715_o;
  wire [23:0] n11716_o;
  wire [24:0] n11717_o;
  wire [24:0] n11718_o;
  wire [23:0] n11719_o;
  wire [23:0] n11720_o;
  wire [24:0] n11721_o;
  wire [24:0] n11722_o;
  wire [23:0] n11723_o;
  wire [23:0] n11724_o;
  wire [24:0] n11725_o;
  wire [24:0] n11726_o;
  wire [23:0] n11727_o;
  wire [23:0] n11728_o;
  wire [24:0] n11729_o;
  wire [24:0] n11730_o;
  wire [24:0] n11731_o;
  wire [24:0] n11732_o;
  wire [24:0] n11733_o;
  wire [2:0] n11734_o;
  wire [24:0] n11735_o;
  wire [31:0] n11736_o;
  wire [23:0] n11737_o;
  wire [23:0] n11738_o;
  wire n11739_o;
  wire [1:0] n11740_o;
  wire n11741_o;
  wire [23:0] n11742_o;
  wire [5:0] n11743_o;
  wire [15:0] n11744_o;
  wire n11745_o;
  wire [1:0] n11746_o;
  wire [1:0] n11747_o;
  wire [23:0] n11748_o;
  wire [23:0] n11749_o;
  wire [23:0] n11750_o;
  wire [23:0] n11751_o;
  wire [24:0] n11752_o;
  wire [24:0] n11753_o;
  wire [23:0] n11754_o;
  wire [23:0] n11755_o;
  wire [24:0] n11756_o;
  wire [24:0] n11757_o;
  wire [23:0] n11758_o;
  wire [23:0] n11759_o;
  wire [24:0] n11760_o;
  wire [24:0] n11761_o;
  wire [23:0] n11762_o;
  wire [23:0] n11763_o;
  wire [24:0] n11764_o;
  wire [24:0] n11765_o;
  wire [23:0] n11766_o;
  wire [23:0] n11767_o;
  wire [24:0] n11768_o;
  wire [24:0] n11769_o;
  wire [24:0] n11770_o;
  wire [24:0] n11771_o;
  wire [24:0] n11772_o;
  wire [2:0] n11773_o;
  wire [24:0] n11774_o;
  wire [31:0] n11775_o;
  wire [23:0] n11776_o;
  wire [23:0] n11777_o;
  wire n11778_o;
  wire [1:0] n11779_o;
  wire n11780_o;
  wire [23:0] n11781_o;
  wire [5:0] n11782_o;
  wire [15:0] n11783_o;
  wire n11784_o;
  wire [1:0] n11785_o;
  wire [1:0] n11786_o;
  wire [23:0] n11787_o;
  wire [23:0] n11788_o;
  wire [1:0] n11856_o;
  assign ready_out = ready;
  assign log1_out = dp_gen_primary_i_n11346;
  assign log1_valid_out = dp_gen_primary_i_n11347;
  assign log2_out = dp_gen_secondary_i_n11630;
  assign log2_valid_out = dp_gen_secondary_i_n11631;
  assign gen_pcore_src_valid_out = n11178_o;
  assign gen_pcore_vm_out = n11179_o;
  assign gen_pcore_fork_out = n11180_o;
  assign gen_pcore_data_flow_out = n11181_o;
  assign gen_pcore_src_stream_out = n11182_o;
  assign gen_pcore_dest_stream_out = n11183_o;
  assign gen_pcore_stream_id_out = n11184_o;
  assign gen_pcore_src_vector_out = n11185_o;
  assign gen_pcore_dst_vector_out = n11186_o;
  assign gen_pcore_src_scatter_out = n11187_o;
  assign gen_pcore_dst_scatter_out = n11188_o;
  assign gen_pcore_src_start_out = n11189_o;
  assign gen_pcore_src_end_out = n11190_o;
  assign gen_pcore_dst_end_out = n11191_o;
  assign gen_pcore_src_addr_out = n11192_o;
  assign gen_pcore_src_addr_mode_out = n11193_o;
  assign gen_pcore_dst_addr_out = n11194_o;
  assign gen_pcore_dst_addr_mode_out = n11195_o;
  assign gen_pcore_src_eof_out = n11196_o;
  assign gen_pcore_bus_id_source_out = n11197_o;
  assign gen_pcore_data_type_source_out = n11198_o;
  assign gen_pcore_data_model_source_out = n11199_o;
  assign gen_pcore_bus_id_dest_out = n11200_o;
  assign gen_pcore_busy_dest_out = n11201_o;
  assign gen_pcore_data_type_dest_out = n11202_o;
  assign gen_pcore_data_model_dest_out = n11203_o;
  assign gen_pcore_src_burstlen_out = n11204_o;
  assign gen_pcore_dst_burstlen_out = n11205_o;
  assign gen_pcore_thread_out = n11206_o;
  assign gen_pcore_mcast_out = n11207_o;
  assign gen_pcore_data_out = n11208_o;
  assign gen_sram_src_valid_out = n11216_o;
  assign gen_sram_vm_out = n11217_o;
  assign gen_sram_fork_out = n11218_o;
  assign gen_sram_data_flow_out = n11219_o;
  assign gen_sram_src_stream_out = n11220_o;
  assign gen_sram_dest_stream_out = n11221_o;
  assign gen_sram_stream_id_out = n11222_o;
  assign gen_sram_src_vector_out = n11223_o;
  assign gen_sram_dst_vector_out = n11224_o;
  assign gen_sram_src_scatter_out = n11225_o;
  assign gen_sram_dst_scatter_out = n11226_o;
  assign gen_sram_src_start_out = n11227_o;
  assign gen_sram_src_end_out = n11228_o;
  assign gen_sram_dst_end_out = n11229_o;
  assign gen_sram_src_addr_out = n11230_o;
  assign gen_sram_src_addr_mode_out = n11231_o;
  assign gen_sram_dst_addr_out = n11232_o;
  assign gen_sram_dst_addr_mode_out = n11233_o;
  assign gen_sram_src_eof_out = n11234_o;
  assign gen_sram_bus_id_source_out = n11235_o;
  assign gen_sram_data_type_source_out = n11236_o;
  assign gen_sram_data_model_source_out = n11237_o;
  assign gen_sram_bus_id_dest_out = n11238_o;
  assign gen_sram_busy_dest_out = n11239_o;
  assign gen_sram_data_type_dest_out = n11240_o;
  assign gen_sram_data_model_dest_out = n11241_o;
  assign gen_sram_src_burstlen_out = n11242_o;
  assign gen_sram_dst_burstlen_out = n11243_o;
  assign gen_sram_thread_out = n11244_o;
  assign gen_sram_mcast_out = n11245_o;
  assign gen_sram_data_out = n11246_o;
  assign gen_ddr_src_valid_out = n11255_o;
  assign gen_ddr_vm_out = n11256_o;
  assign gen_ddr_fork_out = n11257_o;
  assign gen_ddr_data_flow_out = n11258_o;
  assign gen_ddr_src_stream_out = n11259_o;
  assign gen_ddr_dest_stream_out = n11260_o;
  assign gen_ddr_stream_id_out = n11261_o;
  assign gen_ddr_src_vector_out = n11262_o;
  assign gen_ddr_dst_vector_out = n11263_o;
  assign gen_ddr_src_scatter_out = n11264_o;
  assign gen_ddr_dst_scatter_out = n11265_o;
  assign gen_ddr_src_start_out = n11266_o;
  assign gen_ddr_src_end_out = n11267_o;
  assign gen_ddr_dst_end_out = n11268_o;
  assign gen_ddr_src_addr_out = n11269_o;
  assign gen_ddr_src_addr_mode_out = n11270_o;
  assign gen_ddr_dst_addr_out = n11271_o;
  assign gen_ddr_dst_addr_mode_out = n11272_o;
  assign gen_ddr_src_eof_out = n11273_o;
  assign gen_ddr_bus_id_source_out = n11274_o;
  assign gen_ddr_data_type_source_out = n11275_o;
  assign gen_ddr_data_model_source_out = n11276_o;
  assign gen_ddr_bus_id_dest_out = n11277_o;
  assign gen_ddr_busy_dest_out = n11278_o;
  assign gen_ddr_data_type_dest_out = n11279_o;
  assign gen_ddr_data_model_dest_out = n11280_o;
  assign gen_ddr_src_burstlen_out = n11281_o;
  assign gen_ddr_dst_burstlen_out = n11282_o;
  assign gen_ddr_thread_out = n11283_o;
  assign gen_ddr_mcast_out = n11284_o;
  assign gen_ddr_data_out = n11285_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1678:48  */
  assign n11072_o = {instruction_in_stream_process_id, instruction_in_stream_process, instruction_in_dest_addr_mode, instruction_in_source_addr_mode, instruction_in_repeat, instruction_in_data, instruction_in_count, instruction_in_mcast, instruction_in_dest_data_type, instruction_in_dest_bus_id, instruction_in_dest, instruction_in_source_data_type, instruction_in_source_bus_id, instruction_in_source, instruction_in_vm, instruction_in_condition, instruction_in_opcode};
  /* ../../HW/src/dp/dp_fetch.vhd:2156:1  */
  assign n11073_o = {pre_instruction_in_stream_process_id, pre_instruction_in_stream_process, pre_instruction_in_dest_addr_mode, pre_instruction_in_source_addr_mode, pre_instruction_in_repeat, pre_instruction_in_data, pre_instruction_in_count, pre_instruction_in_mcast, pre_instruction_in_dest_data_type, pre_instruction_in_dest_bus_id, pre_instruction_in_dest, pre_instruction_in_source_data_type, pre_instruction_in_source_bus_id, pre_instruction_in_source, pre_instruction_in_vm, pre_instruction_in_condition, pre_instruction_in_opcode};
  /* ../../HW/src/dp/dp_gen_core.vhd:156:8  */
  assign gen_src_valid_1 = dp_gen_primary_i_n11315; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:157:8  */
  assign gen_fork_1 = dp_gen_primary_i_n11317; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:158:8  */
  assign gen_vm_1 = dp_gen_primary_i_n11316; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:159:8  */
  assign gen_data_flow_1 = dp_gen_primary_i_n11318; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:160:8  */
  assign gen_src_stream_1 = dp_gen_primary_i_n11319; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:161:8  */
  assign gen_dest_stream_1 = dp_gen_primary_i_n11320; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:162:8  */
  assign gen_stream_id_1 = dp_gen_primary_i_n11321; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:163:8  */
  assign gen_src_vector_1 = dp_gen_primary_i_n11322; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:164:8  */
  assign gen_dst_vector_1 = dp_gen_primary_i_n11323; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:165:8  */
  assign gen_src_scatter_1 = dp_gen_primary_i_n11324; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:166:8  */
  assign gen_dst_scatter_1 = dp_gen_primary_i_n11325; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:167:8  */
  assign gen_src_start_1 = dp_gen_primary_i_n11326; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:168:8  */
  assign gen_src_end_1 = dp_gen_primary_i_n11327; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:169:8  */
  assign gen_dst_end_1 = dp_gen_primary_i_n11328; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:170:8  */
  assign gen_src_addr_1 = dp_gen_primary_i_n11329; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:171:8  */
  assign gen_src_addr_mode_1 = dp_gen_primary_i_n11330; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:172:8  */
  assign gen_dst_addr_1 = dp_gen_primary_i_n11331; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:173:8  */
  assign gen_dst_addr_mode_1 = dp_gen_primary_i_n11332; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:174:8  */
  assign gen_src_eof_1 = dp_gen_primary_i_n11333; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:175:8  */
  assign gen_bus_id_source_1 = dp_gen_primary_i_n11334; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:176:8  */
  assign gen_data_type_source_1 = dp_gen_primary_i_n11335; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:177:8  */
  assign gen_data_model_source_1 = dp_gen_primary_i_n11336; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:178:8  */
  assign gen_bus_id_dest_1 = dp_gen_primary_i_n11337; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:179:8  */
  assign gen_busy_dest_1 = dp_gen_primary_i_n11338; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:180:8  */
  assign gen_data_type_dest_1 = dp_gen_primary_i_n11339; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:181:8  */
  assign gen_data_model_dest_1 = dp_gen_primary_i_n11340; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:182:8  */
  assign gen_src_burstlen_1 = dp_gen_primary_i_n11341; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:183:8  */
  assign gen_dst_burstlen_1 = dp_gen_primary_i_n11342; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:184:8  */
  assign gen_thread_1 = dp_gen_primary_i_n11343; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:185:8  */
  assign gen_mcast_1 = dp_gen_primary_i_n11344; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:186:8  */
  assign gen_data_1 = dp_gen_primary_i_n11345; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:188:8  */
  assign gen_src_valid_2 = dp_gen_secondary_i_n11599; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:189:8  */
  assign gen_vm_2 = dp_gen_secondary_i_n11600; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:190:8  */
  assign gen_fork_2 = dp_gen_secondary_i_n11601; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:191:8  */
  assign gen_data_flow_2 = dp_gen_secondary_i_n11602; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:192:8  */
  assign gen_src_stream_2 = dp_gen_secondary_i_n11603; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:193:8  */
  assign gen_dest_stream_2 = dp_gen_secondary_i_n11604; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:194:8  */
  assign gen_stream_id_2 = dp_gen_secondary_i_n11605; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:195:8  */
  assign gen_src_vector_2 = dp_gen_secondary_i_n11606; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:196:8  */
  assign gen_dst_vector_2 = dp_gen_secondary_i_n11607; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:197:8  */
  assign gen_src_scatter_2 = dp_gen_secondary_i_n11608; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:198:8  */
  assign gen_dst_scatter_2 = dp_gen_secondary_i_n11609; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:199:8  */
  assign gen_src_start_2 = dp_gen_secondary_i_n11610; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:200:8  */
  assign gen_src_end_2 = dp_gen_secondary_i_n11611; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:201:8  */
  assign gen_dst_end_2 = dp_gen_secondary_i_n11612; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:202:8  */
  assign gen_src_addr_2 = dp_gen_secondary_i_n11613; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:203:8  */
  assign gen_src_addr_mode_2 = dp_gen_secondary_i_n11614; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:204:8  */
  assign gen_dst_addr_2 = dp_gen_secondary_i_n11615; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:205:8  */
  assign gen_dst_addr_mode_2 = dp_gen_secondary_i_n11616; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:206:8  */
  assign gen_src_eof_2 = dp_gen_secondary_i_n11617; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:207:8  */
  assign gen_bus_id_source_2 = dp_gen_secondary_i_n11618; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:208:8  */
  assign gen_data_type_source_2 = dp_gen_secondary_i_n11619; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:209:8  */
  assign gen_data_model_source_2 = dp_gen_secondary_i_n11620; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:210:8  */
  assign gen_bus_id_dest_2 = dp_gen_secondary_i_n11621; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:211:8  */
  assign gen_busy_dest_2 = dp_gen_secondary_i_n11622; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:212:8  */
  assign gen_data_type_dest_2 = dp_gen_secondary_i_n11623; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:213:8  */
  assign gen_data_model_dest_2 = dp_gen_secondary_i_n11624; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:214:8  */
  assign gen_src_burstlen_2 = dp_gen_secondary_i_n11625; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:215:8  */
  assign gen_dst_burstlen_2 = dp_gen_secondary_i_n11626; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:216:8  */
  assign gen_thread_2 = dp_gen_secondary_i_n11627; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:217:8  */
  assign gen_mcast_2 = dp_gen_secondary_i_n11628; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:218:8  */
  assign gen_data_2 = dp_gen_secondary_i_n11629; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:224:8  */
  assign ready = n11856_o; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:266:19  */
  assign n11173_o = gen_src_valid_1[0];
  /* ../../HW/src/dp/dp_gen_core.vhd:268:46  */
  assign n11175_o = gen_src_valid_1[0];
  /* ../../HW/src/dp/dp_gen_core.vhd:301:46  */
  assign n11177_o = gen_src_valid_2[0];
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11178_o = n11173_o ? n11175_o : n11177_o;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11179_o = n11173_o ? gen_vm_1 : gen_vm_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11180_o = n11173_o ? gen_fork_1 : gen_fork_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11181_o = n11173_o ? gen_data_flow_1 : gen_data_flow_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11182_o = n11173_o ? gen_src_stream_1 : gen_src_stream_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11183_o = n11173_o ? gen_dest_stream_1 : gen_dest_stream_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11184_o = n11173_o ? gen_stream_id_1 : gen_stream_id_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11185_o = n11173_o ? gen_src_vector_1 : gen_src_vector_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11186_o = n11173_o ? gen_dst_vector_1 : gen_dst_vector_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11187_o = n11173_o ? gen_src_scatter_1 : gen_src_scatter_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11188_o = n11173_o ? gen_dst_scatter_1 : gen_dst_scatter_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11189_o = n11173_o ? gen_src_start_1 : gen_src_start_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11190_o = n11173_o ? gen_src_end_1 : gen_src_end_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11191_o = n11173_o ? gen_dst_end_1 : gen_dst_end_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11192_o = n11173_o ? gen_src_addr_1 : gen_src_addr_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11193_o = n11173_o ? gen_src_addr_mode_1 : gen_src_addr_mode_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11194_o = n11173_o ? gen_dst_addr_1 : gen_dst_addr_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11195_o = n11173_o ? gen_dst_addr_mode_1 : gen_dst_addr_mode_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11196_o = n11173_o ? gen_src_eof_1 : gen_src_eof_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11197_o = n11173_o ? gen_bus_id_source_1 : gen_bus_id_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11198_o = n11173_o ? gen_data_type_source_1 : gen_data_type_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11199_o = n11173_o ? gen_data_model_source_1 : gen_data_model_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11200_o = n11173_o ? gen_bus_id_dest_1 : gen_bus_id_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11201_o = n11173_o ? gen_busy_dest_1 : gen_busy_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11202_o = n11173_o ? gen_data_type_dest_1 : gen_data_type_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11203_o = n11173_o ? gen_data_model_dest_1 : gen_data_model_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11204_o = n11173_o ? gen_src_burstlen_1 : gen_src_burstlen_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11205_o = n11173_o ? gen_dst_burstlen_1 : gen_dst_burstlen_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11206_o = n11173_o ? gen_thread_1 : gen_thread_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11207_o = n11173_o ? gen_mcast_1 : gen_mcast_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:266:1  */
  assign n11208_o = n11173_o ? gen_data_1 : gen_data_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:19  */
  assign n11213_o = gen_src_valid_1[1];
  /* ../../HW/src/dp/dp_gen_core.vhd:373:45  */
  assign n11214_o = gen_src_valid_1[1];
  /* ../../HW/src/dp/dp_gen_core.vhd:405:45  */
  assign n11215_o = gen_src_valid_2[1];
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11216_o = n11213_o ? n11214_o : n11215_o;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11217_o = n11213_o ? gen_vm_1 : gen_vm_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11218_o = n11213_o ? gen_fork_1 : gen_fork_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11219_o = n11213_o ? gen_data_flow_1 : gen_data_flow_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11220_o = n11213_o ? gen_src_stream_1 : gen_src_stream_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11221_o = n11213_o ? gen_dest_stream_1 : gen_dest_stream_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11222_o = n11213_o ? gen_stream_id_1 : gen_stream_id_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11223_o = n11213_o ? gen_src_vector_1 : gen_src_vector_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11224_o = n11213_o ? gen_dst_vector_1 : gen_dst_vector_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11225_o = n11213_o ? gen_src_scatter_1 : gen_src_scatter_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11226_o = n11213_o ? gen_dst_scatter_1 : gen_dst_scatter_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11227_o = n11213_o ? gen_src_start_1 : gen_src_start_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11228_o = n11213_o ? gen_src_end_1 : gen_src_end_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11229_o = n11213_o ? gen_dst_end_1 : gen_dst_end_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11230_o = n11213_o ? gen_src_addr_1 : gen_src_addr_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11231_o = n11213_o ? gen_src_addr_mode_1 : gen_src_addr_mode_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11232_o = n11213_o ? gen_dst_addr_1 : gen_dst_addr_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11233_o = n11213_o ? gen_dst_addr_mode_1 : gen_dst_addr_mode_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11234_o = n11213_o ? gen_src_eof_1 : gen_src_eof_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11235_o = n11213_o ? gen_bus_id_source_1 : gen_bus_id_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11236_o = n11213_o ? gen_data_type_source_1 : gen_data_type_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11237_o = n11213_o ? gen_data_model_source_1 : gen_data_model_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11238_o = n11213_o ? gen_bus_id_dest_1 : gen_bus_id_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11239_o = n11213_o ? gen_busy_dest_1 : gen_busy_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11240_o = n11213_o ? gen_data_type_dest_1 : gen_data_type_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11241_o = n11213_o ? gen_data_model_dest_1 : gen_data_model_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11242_o = n11213_o ? gen_src_burstlen_1 : gen_src_burstlen_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11243_o = n11213_o ? gen_dst_burstlen_1 : gen_dst_burstlen_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11244_o = n11213_o ? gen_thread_1 : gen_thread_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11245_o = n11213_o ? gen_mcast_1 : gen_mcast_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:372:1  */
  assign n11246_o = n11213_o ? gen_data_1 : gen_data_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:19  */
  assign n11250_o = gen_src_valid_1[2];
  /* ../../HW/src/dp/dp_gen_core.vhd:476:44  */
  assign n11252_o = gen_src_valid_1[2];
  /* ../../HW/src/dp/dp_gen_core.vhd:509:44  */
  assign n11254_o = gen_src_valid_2[2];
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11255_o = n11250_o ? n11252_o : n11254_o;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11256_o = n11250_o ? gen_vm_1 : gen_vm_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11257_o = n11250_o ? gen_fork_1 : gen_fork_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11258_o = n11250_o ? gen_data_flow_1 : gen_data_flow_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11259_o = n11250_o ? gen_src_stream_1 : gen_src_stream_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11260_o = n11250_o ? gen_dest_stream_1 : gen_dest_stream_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11261_o = n11250_o ? gen_stream_id_1 : gen_stream_id_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11262_o = n11250_o ? gen_src_vector_1 : gen_src_vector_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11263_o = n11250_o ? gen_dst_vector_1 : gen_dst_vector_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11264_o = n11250_o ? gen_src_scatter_1 : gen_src_scatter_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11265_o = n11250_o ? gen_dst_scatter_1 : gen_dst_scatter_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11266_o = n11250_o ? gen_src_start_1 : gen_src_start_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11267_o = n11250_o ? gen_src_end_1 : gen_src_end_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11268_o = n11250_o ? gen_dst_end_1 : gen_dst_end_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11269_o = n11250_o ? gen_src_addr_1 : gen_src_addr_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11270_o = n11250_o ? gen_src_addr_mode_1 : gen_src_addr_mode_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11271_o = n11250_o ? gen_dst_addr_1 : gen_dst_addr_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11272_o = n11250_o ? gen_dst_addr_mode_1 : gen_dst_addr_mode_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11273_o = n11250_o ? gen_src_eof_1 : gen_src_eof_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11274_o = n11250_o ? gen_bus_id_source_1 : gen_bus_id_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11275_o = n11250_o ? gen_data_type_source_1 : gen_data_type_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11276_o = n11250_o ? gen_data_model_source_1 : gen_data_model_source_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11277_o = n11250_o ? gen_bus_id_dest_1 : gen_bus_id_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11278_o = n11250_o ? gen_busy_dest_1 : gen_busy_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11279_o = n11250_o ? gen_data_type_dest_1 : gen_data_type_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11280_o = n11250_o ? gen_data_model_dest_1 : gen_data_model_dest_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11281_o = n11250_o ? gen_src_burstlen_1 : gen_src_burstlen_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11282_o = n11250_o ? gen_dst_burstlen_1 : gen_dst_burstlen_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11283_o = n11250_o ? gen_thread_1 : gen_thread_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11284_o = n11250_o ? gen_mcast_1 : gen_mcast_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:474:1  */
  assign n11285_o = n11250_o ? gen_data_1 : gen_data_2;
  /* ../../HW/src/dp/dp_gen_core.vhd:556:40  */
  assign dp_gen_primary_i_n11288 = dp_gen_primary_i_ready_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:557:71  */
  assign n11289_o = instruction_valid_in[0];
  /* ../../HW/src/dp/dp_gen_core.vhd:558:71  */
  assign n11290_o = instruction_valid_in[0];
  /* ../../HW/src/dp/dp_gen_core.vhd:559:67  */
  assign n11291_o = n11072_o[783:8];
  /* ../../HW/src/dp/dp_gen_core.vhd:560:65  */
  assign n11292_o = n11072_o[1563:788];
  /* ../../HW/src/dp/dp_gen_core.vhd:561:75  */
  assign n11293_o = n11072_o[1617];
  /* ../../HW/src/dp/dp_gen_core.vhd:562:78  */
  assign n11294_o = n11072_o[1619:1618];
  /* ../../HW/src/dp/dp_gen_core.vhd:563:63  */
  assign n11295_o = n11072_o[7];
  /* ../../HW/src/dp/dp_gen_core.vhd:564:75  */
  assign n11296_o = n11073_o[783:8];
  /* ../../HW/src/dp/dp_gen_core.vhd:565:73  */
  assign n11297_o = n11073_o[1563:788];
  /* ../../HW/src/dp/dp_gen_core.vhd:566:82  */
  assign n11298_o = n11073_o[785:784];
  /* ../../HW/src/dp/dp_gen_core.vhd:567:80  */
  assign n11299_o = n11073_o[1565:1564];
  /* ../../HW/src/dp/dp_gen_core.vhd:568:77  */
  assign n11300_o = n11072_o[1615];
  /* ../../HW/src/dp/dp_gen_core.vhd:569:75  */
  assign n11301_o = n11072_o[1616];
  /* ../../HW/src/dp/dp_gen_core.vhd:570:74  */
  assign n11302_o = n11072_o[785:784];
  /* ../../HW/src/dp/dp_gen_core.vhd:571:77  */
  assign n11303_o = n11072_o[787:786];
  /* ../../HW/src/dp/dp_gen_core.vhd:572:78  */
  assign n11304_o = n11072_o[783:8];
  /* ../../HW/src/dp/dp_gen_core.vhd:572:85  */
  assign n11305_o = n11304_o[675:674];
  /* ../../HW/src/dp/dp_gen_core.vhd:573:72  */
  assign n11306_o = n11072_o[1565:1564];
  /* ../../HW/src/dp/dp_gen_core.vhd:574:75  */
  assign n11307_o = n11072_o[1567:1566];
  /* ../../HW/src/dp/dp_gen_core.vhd:575:76  */
  assign n11308_o = n11072_o[1563:788];
  /* ../../HW/src/dp/dp_gen_core.vhd:575:81  */
  assign n11309_o = n11308_o[675:674];
  /* ../../HW/src/dp/dp_gen_core.vhd:576:66  */
  assign n11310_o = n11072_o[1573:1568];
  /* ../../HW/src/dp/dp_gen_core.vhd:577:68  */
  assign n11311_o = n11072_o[1597:1574];
  /* ../../HW/src/dp/dp_gen_core.vhd:579:65  */
  assign n11313_o = n11072_o[1613:1598];
  /* ../../HW/src/dp/dp_gen_core.vhd:580:67  */
  assign n11314_o = n11072_o[1614];
  /* ../../HW/src/dp/dp_gen_core.vhd:586:44  */
  assign dp_gen_primary_i_n11315 = dp_gen_primary_i_gen_valid_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:587:41  */
  assign dp_gen_primary_i_n11316 = dp_gen_primary_i_gen_vm_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:588:43  */
  assign dp_gen_primary_i_n11317 = dp_gen_primary_i_gen_fork_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:589:48  */
  assign dp_gen_primary_i_n11318 = dp_gen_primary_i_gen_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:590:49  */
  assign dp_gen_primary_i_n11319 = dp_gen_primary_i_gen_src_stream_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:591:50  */
  assign dp_gen_primary_i_n11320 = dp_gen_primary_i_gen_dest_stream_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:592:50  */
  assign dp_gen_primary_i_n11321 = dp_gen_primary_i_gen_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:593:49  */
  assign dp_gen_primary_i_n11322 = dp_gen_primary_i_gen_src_vector_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:594:49  */
  assign dp_gen_primary_i_n11323 = dp_gen_primary_i_gen_dst_vector_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:595:50  */
  assign dp_gen_primary_i_n11324 = dp_gen_primary_i_gen_src_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:596:50  */
  assign dp_gen_primary_i_n11325 = dp_gen_primary_i_gen_dst_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:597:48  */
  assign dp_gen_primary_i_n11326 = dp_gen_primary_i_gen_src_start_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:598:46  */
  assign dp_gen_primary_i_n11327 = dp_gen_primary_i_gen_src_end_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:599:46  */
  assign dp_gen_primary_i_n11328 = dp_gen_primary_i_gen_dst_end_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:600:50  */
  assign dp_gen_primary_i_n11329 = dp_gen_primary_i_gen_addr_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:601:55  */
  assign dp_gen_primary_i_n11330 = dp_gen_primary_i_gen_addr_source_mode_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:602:48  */
  assign dp_gen_primary_i_n11331 = dp_gen_primary_i_gen_addr_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:603:53  */
  assign dp_gen_primary_i_n11332 = dp_gen_primary_i_gen_addr_dest_mode_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:604:42  */
  assign dp_gen_primary_i_n11333 = dp_gen_primary_i_gen_eof_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:605:52  */
  assign dp_gen_primary_i_n11334 = dp_gen_primary_i_gen_bus_id_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:606:55  */
  assign dp_gen_primary_i_n11335 = dp_gen_primary_i_gen_data_type_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:607:56  */
  assign dp_gen_primary_i_n11336 = dp_gen_primary_i_gen_data_model_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:608:50  */
  assign dp_gen_primary_i_n11337 = dp_gen_primary_i_gen_bus_id_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:609:48  */
  assign dp_gen_primary_i_n11338 = dp_gen_primary_i_gen_busy_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:610:53  */
  assign dp_gen_primary_i_n11339 = dp_gen_primary_i_gen_data_type_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:611:54  */
  assign dp_gen_primary_i_n11340 = dp_gen_primary_i_gen_data_model_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:612:54  */
  assign dp_gen_primary_i_n11341 = dp_gen_primary_i_gen_burstlen_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:613:52  */
  assign dp_gen_primary_i_n11342 = dp_gen_primary_i_gen_burstlen_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:614:45  */
  assign dp_gen_primary_i_n11343 = dp_gen_primary_i_gen_thread_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:615:44  */
  assign dp_gen_primary_i_n11344 = dp_gen_primary_i_gen_mcast_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:616:43  */
  assign dp_gen_primary_i_n11345 = dp_gen_primary_i_gen_data_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:620:38  */
  assign dp_gen_primary_i_n11346 = dp_gen_primary_i_log_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:621:44  */
  assign dp_gen_primary_i_n11347 = dp_gen_primary_i_log_valid_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:546:1  */
  dp_gen_3_0_5b55ec37559bb110228a6591713076b7fa2ce5e8 dp_gen_primary_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_valid_in(n11289_o),
    .instruction_latch_in(n11290_o),
    .instruction_source_in_stride0(n11349_o),
    .instruction_source_in_stride0_count(n11350_o),
    .instruction_source_in_stride0_max(n11351_o),
    .instruction_source_in_stride0_min(n11352_o),
    .instruction_source_in_stride1(n11353_o),
    .instruction_source_in_stride1_count(n11354_o),
    .instruction_source_in_stride1_max(n11355_o),
    .instruction_source_in_stride1_min(n11356_o),
    .instruction_source_in_stride2(n11357_o),
    .instruction_source_in_stride2_count(n11358_o),
    .instruction_source_in_stride2_max(n11359_o),
    .instruction_source_in_stride2_min(n11360_o),
    .instruction_source_in_stride3(n11361_o),
    .instruction_source_in_stride3_count(n11362_o),
    .instruction_source_in_stride3_max(n11363_o),
    .instruction_source_in_stride3_min(n11364_o),
    .instruction_source_in_stride4(n11365_o),
    .instruction_source_in_stride4_count(n11366_o),
    .instruction_source_in_stride4_max(n11367_o),
    .instruction_source_in_stride4_min(n11368_o),
    .instruction_source_in_burst_max(n11369_o),
    .instruction_source_in_burst_max2(n11370_o),
    .instruction_source_in_burst_max_init(n11371_o),
    .instruction_source_in_burst_max_index(n11372_o),
    .instruction_source_in_burst_min(n11373_o),
    .instruction_source_in_bar(n11374_o),
    .instruction_source_in_count(n11375_o),
    .instruction_source_in_burststride(n11376_o),
    .instruction_source_in_double_precision(n11377_o),
    .instruction_source_in_data_model(n11378_o),
    .instruction_source_in_scatter(n11379_o),
    .instruction_source_in_totalcount(n11380_o),
    .instruction_source_in_mcast(n11381_o),
    .instruction_source_in_data(n11382_o),
    .instruction_source_in_repeat(n11383_o),
    .instruction_source_in_datatype(n11384_o),
    .instruction_source_in_bus_id(n11385_o),
    .instruction_source_in_bufsize(n11386_o),
    .instruction_source_in_burst_max_len(n11387_o),
    .instruction_dest_in_stride0(n11388_o),
    .instruction_dest_in_stride0_count(n11389_o),
    .instruction_dest_in_stride0_max(n11390_o),
    .instruction_dest_in_stride0_min(n11391_o),
    .instruction_dest_in_stride1(n11392_o),
    .instruction_dest_in_stride1_count(n11393_o),
    .instruction_dest_in_stride1_max(n11394_o),
    .instruction_dest_in_stride1_min(n11395_o),
    .instruction_dest_in_stride2(n11396_o),
    .instruction_dest_in_stride2_count(n11397_o),
    .instruction_dest_in_stride2_max(n11398_o),
    .instruction_dest_in_stride2_min(n11399_o),
    .instruction_dest_in_stride3(n11400_o),
    .instruction_dest_in_stride3_count(n11401_o),
    .instruction_dest_in_stride3_max(n11402_o),
    .instruction_dest_in_stride3_min(n11403_o),
    .instruction_dest_in_stride4(n11404_o),
    .instruction_dest_in_stride4_count(n11405_o),
    .instruction_dest_in_stride4_max(n11406_o),
    .instruction_dest_in_stride4_min(n11407_o),
    .instruction_dest_in_burst_max(n11408_o),
    .instruction_dest_in_burst_max2(n11409_o),
    .instruction_dest_in_burst_max_init(n11410_o),
    .instruction_dest_in_burst_max_index(n11411_o),
    .instruction_dest_in_burst_min(n11412_o),
    .instruction_dest_in_bar(n11413_o),
    .instruction_dest_in_count(n11414_o),
    .instruction_dest_in_burststride(n11415_o),
    .instruction_dest_in_double_precision(n11416_o),
    .instruction_dest_in_data_model(n11417_o),
    .instruction_dest_in_scatter(n11418_o),
    .instruction_dest_in_totalcount(n11419_o),
    .instruction_dest_in_mcast(n11420_o),
    .instruction_dest_in_data(n11421_o),
    .instruction_dest_in_repeat(n11422_o),
    .instruction_dest_in_datatype(n11423_o),
    .instruction_dest_in_bus_id(n11424_o),
    .instruction_dest_in_bufsize(n11425_o),
    .instruction_dest_in_burst_max_len(n11426_o),
    .instruction_stream_process_in(n11293_o),
    .instruction_stream_process_id_in(n11294_o),
    .instruction_vm_in(n11295_o),
    .pre_instruction_source_in_stride0(n11427_o),
    .pre_instruction_source_in_stride0_count(n11428_o),
    .pre_instruction_source_in_stride0_max(n11429_o),
    .pre_instruction_source_in_stride0_min(n11430_o),
    .pre_instruction_source_in_stride1(n11431_o),
    .pre_instruction_source_in_stride1_count(n11432_o),
    .pre_instruction_source_in_stride1_max(n11433_o),
    .pre_instruction_source_in_stride1_min(n11434_o),
    .pre_instruction_source_in_stride2(n11435_o),
    .pre_instruction_source_in_stride2_count(n11436_o),
    .pre_instruction_source_in_stride2_max(n11437_o),
    .pre_instruction_source_in_stride2_min(n11438_o),
    .pre_instruction_source_in_stride3(n11439_o),
    .pre_instruction_source_in_stride3_count(n11440_o),
    .pre_instruction_source_in_stride3_max(n11441_o),
    .pre_instruction_source_in_stride3_min(n11442_o),
    .pre_instruction_source_in_stride4(n11443_o),
    .pre_instruction_source_in_stride4_count(n11444_o),
    .pre_instruction_source_in_stride4_max(n11445_o),
    .pre_instruction_source_in_stride4_min(n11446_o),
    .pre_instruction_source_in_burst_max(n11447_o),
    .pre_instruction_source_in_burst_max2(n11448_o),
    .pre_instruction_source_in_burst_max_init(n11449_o),
    .pre_instruction_source_in_burst_max_index(n11450_o),
    .pre_instruction_source_in_burst_min(n11451_o),
    .pre_instruction_source_in_bar(n11452_o),
    .pre_instruction_source_in_count(n11453_o),
    .pre_instruction_source_in_burststride(n11454_o),
    .pre_instruction_source_in_double_precision(n11455_o),
    .pre_instruction_source_in_data_model(n11456_o),
    .pre_instruction_source_in_scatter(n11457_o),
    .pre_instruction_source_in_totalcount(n11458_o),
    .pre_instruction_source_in_mcast(n11459_o),
    .pre_instruction_source_in_data(n11460_o),
    .pre_instruction_source_in_repeat(n11461_o),
    .pre_instruction_source_in_datatype(n11462_o),
    .pre_instruction_source_in_bus_id(n11463_o),
    .pre_instruction_source_in_bufsize(n11464_o),
    .pre_instruction_source_in_burst_max_len(n11465_o),
    .pre_instruction_dest_in_stride0(n11466_o),
    .pre_instruction_dest_in_stride0_count(n11467_o),
    .pre_instruction_dest_in_stride0_max(n11468_o),
    .pre_instruction_dest_in_stride0_min(n11469_o),
    .pre_instruction_dest_in_stride1(n11470_o),
    .pre_instruction_dest_in_stride1_count(n11471_o),
    .pre_instruction_dest_in_stride1_max(n11472_o),
    .pre_instruction_dest_in_stride1_min(n11473_o),
    .pre_instruction_dest_in_stride2(n11474_o),
    .pre_instruction_dest_in_stride2_count(n11475_o),
    .pre_instruction_dest_in_stride2_max(n11476_o),
    .pre_instruction_dest_in_stride2_min(n11477_o),
    .pre_instruction_dest_in_stride3(n11478_o),
    .pre_instruction_dest_in_stride3_count(n11479_o),
    .pre_instruction_dest_in_stride3_max(n11480_o),
    .pre_instruction_dest_in_stride3_min(n11481_o),
    .pre_instruction_dest_in_stride4(n11482_o),
    .pre_instruction_dest_in_stride4_count(n11483_o),
    .pre_instruction_dest_in_stride4_max(n11484_o),
    .pre_instruction_dest_in_stride4_min(n11485_o),
    .pre_instruction_dest_in_burst_max(n11486_o),
    .pre_instruction_dest_in_burst_max2(n11487_o),
    .pre_instruction_dest_in_burst_max_init(n11488_o),
    .pre_instruction_dest_in_burst_max_index(n11489_o),
    .pre_instruction_dest_in_burst_min(n11490_o),
    .pre_instruction_dest_in_bar(n11491_o),
    .pre_instruction_dest_in_count(n11492_o),
    .pre_instruction_dest_in_burststride(n11493_o),
    .pre_instruction_dest_in_double_precision(n11494_o),
    .pre_instruction_dest_in_data_model(n11495_o),
    .pre_instruction_dest_in_scatter(n11496_o),
    .pre_instruction_dest_in_totalcount(n11497_o),
    .pre_instruction_dest_in_mcast(n11498_o),
    .pre_instruction_dest_in_data(n11499_o),
    .pre_instruction_dest_in_repeat(n11500_o),
    .pre_instruction_dest_in_datatype(n11501_o),
    .pre_instruction_dest_in_bus_id(n11502_o),
    .pre_instruction_dest_in_bufsize(n11503_o),
    .pre_instruction_dest_in_burst_max_len(n11504_o),
    .pre_instruction_bus_id_source_in(n11298_o),
    .pre_instruction_bus_id_dest_in(n11299_o),
    .instruction_source_addr_mode_in(n11300_o),
    .instruction_dest_addr_mode_in(n11301_o),
    .instruction_bus_id_source_in(n11302_o),
    .instruction_data_type_source_in(n11303_o),
    .instruction_data_model_source_in(n11305_o),
    .instruction_bus_id_dest_in(n11306_o),
    .instruction_data_type_dest_in(n11307_o),
    .instruction_data_model_dest_in(n11309_o),
    .instruction_gen_len_in(n11311_o),
    .instruction_mcast_in(n11310_o),
    .instruction_thread_in(n11312_o),
    .instruction_data_in(n11313_o),
    .instruction_repeat_in(n11314_o),
    .wr_maxburstlen_in(wr_maxburstlen_in),
    .wr_full_in(full_in),
    .waitreq_in(waitreq_in),
    .gen_bar_in(bar_in),
    .ready_out(dp_gen_primary_i_ready_out),
    .gen_valid_out(dp_gen_primary_i_gen_valid_out),
    .gen_vm_out(dp_gen_primary_i_gen_vm_out),
    .gen_fork_out(dp_gen_primary_i_gen_fork_out),
    .gen_data_flow_out(dp_gen_primary_i_gen_data_flow_out),
    .gen_src_stream_out(dp_gen_primary_i_gen_src_stream_out),
    .gen_dest_stream_out(dp_gen_primary_i_gen_dest_stream_out),
    .gen_stream_id_out(dp_gen_primary_i_gen_stream_id_out),
    .gen_src_vector_out(dp_gen_primary_i_gen_src_vector_out),
    .gen_dst_vector_out(dp_gen_primary_i_gen_dst_vector_out),
    .gen_src_scatter_out(dp_gen_primary_i_gen_src_scatter_out),
    .gen_dst_scatter_out(dp_gen_primary_i_gen_dst_scatter_out),
    .gen_src_start_out(dp_gen_primary_i_gen_src_start_out),
    .gen_src_end_out(dp_gen_primary_i_gen_src_end_out),
    .gen_dst_end_out(dp_gen_primary_i_gen_dst_end_out),
    .gen_addr_source_out(dp_gen_primary_i_gen_addr_source_out),
    .gen_addr_source_mode_out(dp_gen_primary_i_gen_addr_source_mode_out),
    .gen_addr_dest_out(dp_gen_primary_i_gen_addr_dest_out),
    .gen_addr_dest_mode_out(dp_gen_primary_i_gen_addr_dest_mode_out),
    .gen_eof_out(dp_gen_primary_i_gen_eof_out),
    .gen_bus_id_source_out(dp_gen_primary_i_gen_bus_id_source_out),
    .gen_data_type_source_out(dp_gen_primary_i_gen_data_type_source_out),
    .gen_data_model_source_out(dp_gen_primary_i_gen_data_model_source_out),
    .gen_bus_id_dest_out(dp_gen_primary_i_gen_bus_id_dest_out),
    .gen_busy_dest_out(dp_gen_primary_i_gen_busy_dest_out),
    .gen_data_type_dest_out(dp_gen_primary_i_gen_data_type_dest_out),
    .gen_data_model_dest_out(dp_gen_primary_i_gen_data_model_dest_out),
    .gen_burstlen_source_out(dp_gen_primary_i_gen_burstlen_source_out),
    .gen_burstlen_dest_out(dp_gen_primary_i_gen_burstlen_dest_out),
    .gen_thread_out(dp_gen_primary_i_gen_thread_out),
    .gen_mcast_out(dp_gen_primary_i_gen_mcast_out),
    .gen_data_out(dp_gen_primary_i_gen_data_out),
    .log_out(dp_gen_primary_i_log_out),
    .log_valid_out(dp_gen_primary_i_log_valid_out));
  assign n11349_o = n11291_o[23:0];
  assign n11350_o = n11291_o[47:24];
  assign n11351_o = n11291_o[72:48];
  assign n11352_o = n11291_o[97:73];
  assign n11353_o = n11291_o[121:98];
  assign n11354_o = n11291_o[145:122];
  assign n11355_o = n11291_o[170:146];
  assign n11356_o = n11291_o[195:171];
  assign n11357_o = n11291_o[219:196];
  assign n11358_o = n11291_o[243:220];
  assign n11359_o = n11291_o[268:244];
  assign n11360_o = n11291_o[293:269];
  assign n11361_o = n11291_o[317:294];
  assign n11362_o = n11291_o[341:318];
  assign n11363_o = n11291_o[366:342];
  assign n11364_o = n11291_o[391:367];
  assign n11365_o = n11291_o[415:392];
  assign n11366_o = n11291_o[439:416];
  assign n11367_o = n11291_o[464:440];
  assign n11368_o = n11291_o[489:465];
  assign n11369_o = n11291_o[514:490];
  assign n11370_o = n11291_o[539:515];
  assign n11371_o = n11291_o[564:540];
  assign n11372_o = n11291_o[567:565];
  assign n11373_o = n11291_o[592:568];
  assign n11374_o = n11291_o[624:593];
  assign n11375_o = n11291_o[648:625];
  assign n11376_o = n11291_o[672:649];
  assign n11377_o = n11291_o[673];
  assign n11378_o = n11291_o[675:674];
  assign n11379_o = n11291_o[676];
  assign n11380_o = n11291_o[700:677];
  assign n11381_o = n11291_o[706:701];
  assign n11382_o = n11291_o[722:707];
  assign n11383_o = n11291_o[723];
  assign n11384_o = n11291_o[725:724];
  assign n11385_o = n11291_o[727:726];
  assign n11386_o = n11291_o[751:728];
  assign n11387_o = n11291_o[775:752];
  assign n11388_o = n11292_o[23:0];
  assign n11389_o = n11292_o[47:24];
  assign n11390_o = n11292_o[72:48];
  assign n11391_o = n11292_o[97:73];
  assign n11392_o = n11292_o[121:98];
  assign n11393_o = n11292_o[145:122];
  assign n11394_o = n11292_o[170:146];
  assign n11395_o = n11292_o[195:171];
  assign n11396_o = n11292_o[219:196];
  assign n11397_o = n11292_o[243:220];
  assign n11398_o = n11292_o[268:244];
  assign n11399_o = n11292_o[293:269];
  assign n11400_o = n11292_o[317:294];
  assign n11401_o = n11292_o[341:318];
  assign n11402_o = n11292_o[366:342];
  assign n11403_o = n11292_o[391:367];
  assign n11404_o = n11292_o[415:392];
  assign n11405_o = n11292_o[439:416];
  assign n11406_o = n11292_o[464:440];
  assign n11407_o = n11292_o[489:465];
  assign n11408_o = n11292_o[514:490];
  assign n11409_o = n11292_o[539:515];
  assign n11410_o = n11292_o[564:540];
  /* ../../HW/src/dp/dp_fetch.vhd:612:10  */
  assign n11411_o = n11292_o[567:565];
  assign n11412_o = n11292_o[592:568];
  /* ../../HW/src/dp/dp_fetch.vhd:611:10  */
  assign n11413_o = n11292_o[624:593];
  assign n11414_o = n11292_o[648:625];
  /* ../../HW/src/dp/dp_fetch.vhd:610:10  */
  assign n11415_o = n11292_o[672:649];
  /* ../../HW/src/dp/dp_fetch.vhd:610:10  */
  assign n11416_o = n11292_o[673];
  assign n11417_o = n11292_o[675:674];
  /* ../../HW/src/dp/dp_fetch.vhd:610:10  */
  assign n11418_o = n11292_o[676];
  assign n11419_o = n11292_o[700:677];
  /* ../../HW/src/dp/dp_fetch.vhd:786:10  */
  assign n11420_o = n11292_o[706:701];
  assign n11421_o = n11292_o[722:707];
  /* ../../HW/src/dp/dp_fetch.vhd:785:10  */
  assign n11422_o = n11292_o[723];
  assign n11423_o = n11292_o[725:724];
  /* ../../HW/src/dp/dp_fetch.vhd:784:10  */
  assign n11424_o = n11292_o[727:726];
  /* ../../HW/src/dp/dp_fetch.vhd:784:10  */
  assign n11425_o = n11292_o[751:728];
  assign n11426_o = n11292_o[775:752];
  /* ../../HW/src/dp/dp_fetch.vhd:784:10  */
  assign n11427_o = n11296_o[23:0];
  assign n11428_o = n11296_o[47:24];
  assign n11429_o = n11296_o[72:48];
  assign n11430_o = n11296_o[97:73];
  assign n11431_o = n11296_o[121:98];
  assign n11432_o = n11296_o[145:122];
  assign n11433_o = n11296_o[170:146];
  assign n11434_o = n11296_o[195:171];
  assign n11435_o = n11296_o[219:196];
  assign n11436_o = n11296_o[243:220];
  assign n11437_o = n11296_o[268:244];
  assign n11438_o = n11296_o[293:269];
  assign n11439_o = n11296_o[317:294];
  assign n11440_o = n11296_o[341:318];
  assign n11441_o = n11296_o[366:342];
  assign n11442_o = n11296_o[391:367];
  assign n11443_o = n11296_o[415:392];
  assign n11444_o = n11296_o[439:416];
  assign n11445_o = n11296_o[464:440];
  assign n11446_o = n11296_o[489:465];
  assign n11447_o = n11296_o[514:490];
  assign n11448_o = n11296_o[539:515];
  assign n11449_o = n11296_o[564:540];
  assign n11450_o = n11296_o[567:565];
  assign n11451_o = n11296_o[592:568];
  assign n11452_o = n11296_o[624:593];
  assign n11453_o = n11296_o[648:625];
  assign n11454_o = n11296_o[672:649];
  assign n11455_o = n11296_o[673];
  assign n11456_o = n11296_o[675:674];
  assign n11457_o = n11296_o[676];
  assign n11458_o = n11296_o[700:677];
  assign n11459_o = n11296_o[706:701];
  assign n11460_o = n11296_o[722:707];
  assign n11461_o = n11296_o[723];
  assign n11462_o = n11296_o[725:724];
  assign n11463_o = n11296_o[727:726];
  assign n11464_o = n11296_o[751:728];
  assign n11465_o = n11296_o[775:752];
  assign n11466_o = n11297_o[23:0];
  assign n11467_o = n11297_o[47:24];
  assign n11468_o = n11297_o[72:48];
  assign n11469_o = n11297_o[97:73];
  assign n11470_o = n11297_o[121:98];
  assign n11471_o = n11297_o[145:122];
  assign n11472_o = n11297_o[170:146];
  assign n11473_o = n11297_o[195:171];
  assign n11474_o = n11297_o[219:196];
  assign n11475_o = n11297_o[243:220];
  assign n11476_o = n11297_o[268:244];
  assign n11477_o = n11297_o[293:269];
  assign n11478_o = n11297_o[317:294];
  assign n11479_o = n11297_o[341:318];
  assign n11480_o = n11297_o[366:342];
  assign n11481_o = n11297_o[391:367];
  assign n11482_o = n11297_o[415:392];
  assign n11483_o = n11297_o[439:416];
  assign n11484_o = n11297_o[464:440];
  assign n11485_o = n11297_o[489:465];
  assign n11486_o = n11297_o[514:490];
  assign n11487_o = n11297_o[539:515];
  assign n11488_o = n11297_o[564:540];
  assign n11489_o = n11297_o[567:565];
  assign n11490_o = n11297_o[592:568];
  assign n11491_o = n11297_o[624:593];
  assign n11492_o = n11297_o[648:625];
  assign n11493_o = n11297_o[672:649];
  assign n11494_o = n11297_o[673];
  assign n11495_o = n11297_o[675:674];
  assign n11496_o = n11297_o[676];
  assign n11497_o = n11297_o[700:677];
  assign n11498_o = n11297_o[706:701];
  assign n11499_o = n11297_o[722:707];
  assign n11500_o = n11297_o[723];
  assign n11501_o = n11297_o[725:724];
  assign n11502_o = n11297_o[727:726];
  assign n11503_o = n11297_o[751:728];
  assign n11504_o = n11297_o[775:752];
  /* ../../HW/src/dp/dp_gen_core.vhd:634:40  */
  assign dp_gen_secondary_i_n11572 = dp_gen_secondary_i_ready_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:635:71  */
  assign n11573_o = instruction_valid_in[1];
  /* ../../HW/src/dp/dp_gen_core.vhd:636:71  */
  assign n11574_o = instruction_valid_in[1];
  /* ../../HW/src/dp/dp_gen_core.vhd:637:67  */
  assign n11575_o = n11072_o[783:8];
  /* ../../HW/src/dp/dp_gen_core.vhd:638:65  */
  assign n11576_o = n11072_o[1563:788];
  /* ../../HW/src/dp/dp_gen_core.vhd:639:75  */
  assign n11577_o = n11072_o[1617];
  /* ../../HW/src/dp/dp_gen_core.vhd:640:78  */
  assign n11578_o = n11072_o[1619:1618];
  /* ../../HW/src/dp/dp_gen_core.vhd:641:63  */
  assign n11579_o = n11072_o[7];
  /* ../../HW/src/dp/dp_gen_core.vhd:642:75  */
  assign n11580_o = n11073_o[783:8];
  /* ../../HW/src/dp/dp_gen_core.vhd:643:73  */
  assign n11581_o = n11073_o[1563:788];
  /* ../../HW/src/dp/dp_gen_core.vhd:644:82  */
  assign n11582_o = n11073_o[785:784];
  /* ../../HW/src/dp/dp_gen_core.vhd:645:80  */
  assign n11583_o = n11073_o[1565:1564];
  /* ../../HW/src/dp/dp_gen_core.vhd:646:77  */
  assign n11584_o = n11072_o[1615];
  /* ../../HW/src/dp/dp_gen_core.vhd:647:75  */
  assign n11585_o = n11072_o[1616];
  /* ../../HW/src/dp/dp_gen_core.vhd:648:74  */
  assign n11586_o = n11072_o[785:784];
  /* ../../HW/src/dp/dp_gen_core.vhd:649:77  */
  assign n11587_o = n11072_o[787:786];
  /* ../../HW/src/dp/dp_gen_core.vhd:650:78  */
  assign n11588_o = n11072_o[783:8];
  /* ../../HW/src/dp/dp_gen_core.vhd:650:85  */
  assign n11589_o = n11588_o[675:674];
  /* ../../HW/src/dp/dp_gen_core.vhd:651:72  */
  assign n11590_o = n11072_o[1565:1564];
  /* ../../HW/src/dp/dp_gen_core.vhd:652:75  */
  assign n11591_o = n11072_o[1567:1566];
  /* ../../HW/src/dp/dp_gen_core.vhd:653:76  */
  assign n11592_o = n11072_o[1563:788];
  /* ../../HW/src/dp/dp_gen_core.vhd:653:81  */
  assign n11593_o = n11592_o[675:674];
  /* ../../HW/src/dp/dp_gen_core.vhd:654:66  */
  assign n11594_o = n11072_o[1573:1568];
  /* ../../HW/src/dp/dp_gen_core.vhd:655:68  */
  assign n11595_o = n11072_o[1597:1574];
  /* ../../HW/src/dp/dp_gen_core.vhd:657:65  */
  assign n11597_o = n11072_o[1613:1598];
  /* ../../HW/src/dp/dp_gen_core.vhd:658:67  */
  assign n11598_o = n11072_o[1614];
  /* ../../HW/src/dp/dp_gen_core.vhd:665:44  */
  assign dp_gen_secondary_i_n11599 = dp_gen_secondary_i_gen_valid_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:666:41  */
  assign dp_gen_secondary_i_n11600 = dp_gen_secondary_i_gen_vm_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:667:43  */
  assign dp_gen_secondary_i_n11601 = dp_gen_secondary_i_gen_fork_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:668:48  */
  assign dp_gen_secondary_i_n11602 = dp_gen_secondary_i_gen_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:669:49  */
  assign dp_gen_secondary_i_n11603 = dp_gen_secondary_i_gen_src_stream_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:670:50  */
  assign dp_gen_secondary_i_n11604 = dp_gen_secondary_i_gen_dest_stream_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:671:50  */
  assign dp_gen_secondary_i_n11605 = dp_gen_secondary_i_gen_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:672:49  */
  assign dp_gen_secondary_i_n11606 = dp_gen_secondary_i_gen_src_vector_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:673:49  */
  assign dp_gen_secondary_i_n11607 = dp_gen_secondary_i_gen_dst_vector_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:674:50  */
  assign dp_gen_secondary_i_n11608 = dp_gen_secondary_i_gen_src_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:675:50  */
  assign dp_gen_secondary_i_n11609 = dp_gen_secondary_i_gen_dst_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:676:48  */
  assign dp_gen_secondary_i_n11610 = dp_gen_secondary_i_gen_src_start_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:677:46  */
  assign dp_gen_secondary_i_n11611 = dp_gen_secondary_i_gen_src_end_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:678:46  */
  assign dp_gen_secondary_i_n11612 = dp_gen_secondary_i_gen_dst_end_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:679:50  */
  assign dp_gen_secondary_i_n11613 = dp_gen_secondary_i_gen_addr_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:680:55  */
  assign dp_gen_secondary_i_n11614 = dp_gen_secondary_i_gen_addr_source_mode_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:681:48  */
  assign dp_gen_secondary_i_n11615 = dp_gen_secondary_i_gen_addr_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:682:53  */
  assign dp_gen_secondary_i_n11616 = dp_gen_secondary_i_gen_addr_dest_mode_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:683:42  */
  assign dp_gen_secondary_i_n11617 = dp_gen_secondary_i_gen_eof_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:684:52  */
  assign dp_gen_secondary_i_n11618 = dp_gen_secondary_i_gen_bus_id_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:685:55  */
  assign dp_gen_secondary_i_n11619 = dp_gen_secondary_i_gen_data_type_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:686:56  */
  assign dp_gen_secondary_i_n11620 = dp_gen_secondary_i_gen_data_model_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:687:50  */
  assign dp_gen_secondary_i_n11621 = dp_gen_secondary_i_gen_bus_id_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:688:48  */
  assign dp_gen_secondary_i_n11622 = dp_gen_secondary_i_gen_busy_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:689:53  */
  assign dp_gen_secondary_i_n11623 = dp_gen_secondary_i_gen_data_type_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:690:54  */
  assign dp_gen_secondary_i_n11624 = dp_gen_secondary_i_gen_data_model_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:691:54  */
  assign dp_gen_secondary_i_n11625 = dp_gen_secondary_i_gen_burstlen_source_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:692:52  */
  assign dp_gen_secondary_i_n11626 = dp_gen_secondary_i_gen_burstlen_dest_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:693:45  */
  assign dp_gen_secondary_i_n11627 = dp_gen_secondary_i_gen_thread_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:694:44  */
  assign dp_gen_secondary_i_n11628 = dp_gen_secondary_i_gen_mcast_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:695:43  */
  assign dp_gen_secondary_i_n11629 = dp_gen_secondary_i_gen_data_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:699:38  */
  assign dp_gen_secondary_i_n11630 = dp_gen_secondary_i_log_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:700:44  */
  assign dp_gen_secondary_i_n11631 = dp_gen_secondary_i_log_valid_out; // (signal)
  /* ../../HW/src/dp/dp_gen_core.vhd:624:1  */
  dp_gen_3_1_5b55ec37559bb110228a6591713076b7fa2ce5e8 dp_gen_secondary_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_valid_in(n11573_o),
    .instruction_latch_in(n11574_o),
    .instruction_source_in_stride0(n11633_o),
    .instruction_source_in_stride0_count(n11634_o),
    .instruction_source_in_stride0_max(n11635_o),
    .instruction_source_in_stride0_min(n11636_o),
    .instruction_source_in_stride1(n11637_o),
    .instruction_source_in_stride1_count(n11638_o),
    .instruction_source_in_stride1_max(n11639_o),
    .instruction_source_in_stride1_min(n11640_o),
    .instruction_source_in_stride2(n11641_o),
    .instruction_source_in_stride2_count(n11642_o),
    .instruction_source_in_stride2_max(n11643_o),
    .instruction_source_in_stride2_min(n11644_o),
    .instruction_source_in_stride3(n11645_o),
    .instruction_source_in_stride3_count(n11646_o),
    .instruction_source_in_stride3_max(n11647_o),
    .instruction_source_in_stride3_min(n11648_o),
    .instruction_source_in_stride4(n11649_o),
    .instruction_source_in_stride4_count(n11650_o),
    .instruction_source_in_stride4_max(n11651_o),
    .instruction_source_in_stride4_min(n11652_o),
    .instruction_source_in_burst_max(n11653_o),
    .instruction_source_in_burst_max2(n11654_o),
    .instruction_source_in_burst_max_init(n11655_o),
    .instruction_source_in_burst_max_index(n11656_o),
    .instruction_source_in_burst_min(n11657_o),
    .instruction_source_in_bar(n11658_o),
    .instruction_source_in_count(n11659_o),
    .instruction_source_in_burststride(n11660_o),
    .instruction_source_in_double_precision(n11661_o),
    .instruction_source_in_data_model(n11662_o),
    .instruction_source_in_scatter(n11663_o),
    .instruction_source_in_totalcount(n11664_o),
    .instruction_source_in_mcast(n11665_o),
    .instruction_source_in_data(n11666_o),
    .instruction_source_in_repeat(n11667_o),
    .instruction_source_in_datatype(n11668_o),
    .instruction_source_in_bus_id(n11669_o),
    .instruction_source_in_bufsize(n11670_o),
    .instruction_source_in_burst_max_len(n11671_o),
    .instruction_dest_in_stride0(n11672_o),
    .instruction_dest_in_stride0_count(n11673_o),
    .instruction_dest_in_stride0_max(n11674_o),
    .instruction_dest_in_stride0_min(n11675_o),
    .instruction_dest_in_stride1(n11676_o),
    .instruction_dest_in_stride1_count(n11677_o),
    .instruction_dest_in_stride1_max(n11678_o),
    .instruction_dest_in_stride1_min(n11679_o),
    .instruction_dest_in_stride2(n11680_o),
    .instruction_dest_in_stride2_count(n11681_o),
    .instruction_dest_in_stride2_max(n11682_o),
    .instruction_dest_in_stride2_min(n11683_o),
    .instruction_dest_in_stride3(n11684_o),
    .instruction_dest_in_stride3_count(n11685_o),
    .instruction_dest_in_stride3_max(n11686_o),
    .instruction_dest_in_stride3_min(n11687_o),
    .instruction_dest_in_stride4(n11688_o),
    .instruction_dest_in_stride4_count(n11689_o),
    .instruction_dest_in_stride4_max(n11690_o),
    .instruction_dest_in_stride4_min(n11691_o),
    .instruction_dest_in_burst_max(n11692_o),
    .instruction_dest_in_burst_max2(n11693_o),
    .instruction_dest_in_burst_max_init(n11694_o),
    .instruction_dest_in_burst_max_index(n11695_o),
    .instruction_dest_in_burst_min(n11696_o),
    .instruction_dest_in_bar(n11697_o),
    .instruction_dest_in_count(n11698_o),
    .instruction_dest_in_burststride(n11699_o),
    .instruction_dest_in_double_precision(n11700_o),
    .instruction_dest_in_data_model(n11701_o),
    .instruction_dest_in_scatter(n11702_o),
    .instruction_dest_in_totalcount(n11703_o),
    .instruction_dest_in_mcast(n11704_o),
    .instruction_dest_in_data(n11705_o),
    .instruction_dest_in_repeat(n11706_o),
    .instruction_dest_in_datatype(n11707_o),
    .instruction_dest_in_bus_id(n11708_o),
    .instruction_dest_in_bufsize(n11709_o),
    .instruction_dest_in_burst_max_len(n11710_o),
    .instruction_stream_process_in(n11577_o),
    .instruction_stream_process_id_in(n11578_o),
    .instruction_vm_in(n11579_o),
    .pre_instruction_source_in_stride0(n11711_o),
    .pre_instruction_source_in_stride0_count(n11712_o),
    .pre_instruction_source_in_stride0_max(n11713_o),
    .pre_instruction_source_in_stride0_min(n11714_o),
    .pre_instruction_source_in_stride1(n11715_o),
    .pre_instruction_source_in_stride1_count(n11716_o),
    .pre_instruction_source_in_stride1_max(n11717_o),
    .pre_instruction_source_in_stride1_min(n11718_o),
    .pre_instruction_source_in_stride2(n11719_o),
    .pre_instruction_source_in_stride2_count(n11720_o),
    .pre_instruction_source_in_stride2_max(n11721_o),
    .pre_instruction_source_in_stride2_min(n11722_o),
    .pre_instruction_source_in_stride3(n11723_o),
    .pre_instruction_source_in_stride3_count(n11724_o),
    .pre_instruction_source_in_stride3_max(n11725_o),
    .pre_instruction_source_in_stride3_min(n11726_o),
    .pre_instruction_source_in_stride4(n11727_o),
    .pre_instruction_source_in_stride4_count(n11728_o),
    .pre_instruction_source_in_stride4_max(n11729_o),
    .pre_instruction_source_in_stride4_min(n11730_o),
    .pre_instruction_source_in_burst_max(n11731_o),
    .pre_instruction_source_in_burst_max2(n11732_o),
    .pre_instruction_source_in_burst_max_init(n11733_o),
    .pre_instruction_source_in_burst_max_index(n11734_o),
    .pre_instruction_source_in_burst_min(n11735_o),
    .pre_instruction_source_in_bar(n11736_o),
    .pre_instruction_source_in_count(n11737_o),
    .pre_instruction_source_in_burststride(n11738_o),
    .pre_instruction_source_in_double_precision(n11739_o),
    .pre_instruction_source_in_data_model(n11740_o),
    .pre_instruction_source_in_scatter(n11741_o),
    .pre_instruction_source_in_totalcount(n11742_o),
    .pre_instruction_source_in_mcast(n11743_o),
    .pre_instruction_source_in_data(n11744_o),
    .pre_instruction_source_in_repeat(n11745_o),
    .pre_instruction_source_in_datatype(n11746_o),
    .pre_instruction_source_in_bus_id(n11747_o),
    .pre_instruction_source_in_bufsize(n11748_o),
    .pre_instruction_source_in_burst_max_len(n11749_o),
    .pre_instruction_dest_in_stride0(n11750_o),
    .pre_instruction_dest_in_stride0_count(n11751_o),
    .pre_instruction_dest_in_stride0_max(n11752_o),
    .pre_instruction_dest_in_stride0_min(n11753_o),
    .pre_instruction_dest_in_stride1(n11754_o),
    .pre_instruction_dest_in_stride1_count(n11755_o),
    .pre_instruction_dest_in_stride1_max(n11756_o),
    .pre_instruction_dest_in_stride1_min(n11757_o),
    .pre_instruction_dest_in_stride2(n11758_o),
    .pre_instruction_dest_in_stride2_count(n11759_o),
    .pre_instruction_dest_in_stride2_max(n11760_o),
    .pre_instruction_dest_in_stride2_min(n11761_o),
    .pre_instruction_dest_in_stride3(n11762_o),
    .pre_instruction_dest_in_stride3_count(n11763_o),
    .pre_instruction_dest_in_stride3_max(n11764_o),
    .pre_instruction_dest_in_stride3_min(n11765_o),
    .pre_instruction_dest_in_stride4(n11766_o),
    .pre_instruction_dest_in_stride4_count(n11767_o),
    .pre_instruction_dest_in_stride4_max(n11768_o),
    .pre_instruction_dest_in_stride4_min(n11769_o),
    .pre_instruction_dest_in_burst_max(n11770_o),
    .pre_instruction_dest_in_burst_max2(n11771_o),
    .pre_instruction_dest_in_burst_max_init(n11772_o),
    .pre_instruction_dest_in_burst_max_index(n11773_o),
    .pre_instruction_dest_in_burst_min(n11774_o),
    .pre_instruction_dest_in_bar(n11775_o),
    .pre_instruction_dest_in_count(n11776_o),
    .pre_instruction_dest_in_burststride(n11777_o),
    .pre_instruction_dest_in_double_precision(n11778_o),
    .pre_instruction_dest_in_data_model(n11779_o),
    .pre_instruction_dest_in_scatter(n11780_o),
    .pre_instruction_dest_in_totalcount(n11781_o),
    .pre_instruction_dest_in_mcast(n11782_o),
    .pre_instruction_dest_in_data(n11783_o),
    .pre_instruction_dest_in_repeat(n11784_o),
    .pre_instruction_dest_in_datatype(n11785_o),
    .pre_instruction_dest_in_bus_id(n11786_o),
    .pre_instruction_dest_in_bufsize(n11787_o),
    .pre_instruction_dest_in_burst_max_len(n11788_o),
    .pre_instruction_bus_id_source_in(n11582_o),
    .pre_instruction_bus_id_dest_in(n11583_o),
    .instruction_source_addr_mode_in(n11584_o),
    .instruction_dest_addr_mode_in(n11585_o),
    .instruction_bus_id_source_in(n11586_o),
    .instruction_data_type_source_in(n11587_o),
    .instruction_data_model_source_in(n11589_o),
    .instruction_bus_id_dest_in(n11590_o),
    .instruction_data_type_dest_in(n11591_o),
    .instruction_data_model_dest_in(n11593_o),
    .instruction_gen_len_in(n11595_o),
    .instruction_mcast_in(n11594_o),
    .instruction_thread_in(n11596_o),
    .instruction_data_in(n11597_o),
    .instruction_repeat_in(n11598_o),
    .wr_maxburstlen_in(wr_maxburstlen_in),
    .wr_full_in(full_in),
    .waitreq_in(waitreq_in),
    .gen_bar_in(bar_in),
    .ready_out(dp_gen_secondary_i_ready_out),
    .gen_valid_out(dp_gen_secondary_i_gen_valid_out),
    .gen_vm_out(dp_gen_secondary_i_gen_vm_out),
    .gen_fork_out(dp_gen_secondary_i_gen_fork_out),
    .gen_data_flow_out(dp_gen_secondary_i_gen_data_flow_out),
    .gen_src_stream_out(dp_gen_secondary_i_gen_src_stream_out),
    .gen_dest_stream_out(dp_gen_secondary_i_gen_dest_stream_out),
    .gen_stream_id_out(dp_gen_secondary_i_gen_stream_id_out),
    .gen_src_vector_out(dp_gen_secondary_i_gen_src_vector_out),
    .gen_dst_vector_out(dp_gen_secondary_i_gen_dst_vector_out),
    .gen_src_scatter_out(dp_gen_secondary_i_gen_src_scatter_out),
    .gen_dst_scatter_out(dp_gen_secondary_i_gen_dst_scatter_out),
    .gen_src_start_out(dp_gen_secondary_i_gen_src_start_out),
    .gen_src_end_out(dp_gen_secondary_i_gen_src_end_out),
    .gen_dst_end_out(dp_gen_secondary_i_gen_dst_end_out),
    .gen_addr_source_out(dp_gen_secondary_i_gen_addr_source_out),
    .gen_addr_source_mode_out(dp_gen_secondary_i_gen_addr_source_mode_out),
    .gen_addr_dest_out(dp_gen_secondary_i_gen_addr_dest_out),
    .gen_addr_dest_mode_out(dp_gen_secondary_i_gen_addr_dest_mode_out),
    .gen_eof_out(dp_gen_secondary_i_gen_eof_out),
    .gen_bus_id_source_out(dp_gen_secondary_i_gen_bus_id_source_out),
    .gen_data_type_source_out(dp_gen_secondary_i_gen_data_type_source_out),
    .gen_data_model_source_out(dp_gen_secondary_i_gen_data_model_source_out),
    .gen_bus_id_dest_out(dp_gen_secondary_i_gen_bus_id_dest_out),
    .gen_busy_dest_out(dp_gen_secondary_i_gen_busy_dest_out),
    .gen_data_type_dest_out(dp_gen_secondary_i_gen_data_type_dest_out),
    .gen_data_model_dest_out(dp_gen_secondary_i_gen_data_model_dest_out),
    .gen_burstlen_source_out(dp_gen_secondary_i_gen_burstlen_source_out),
    .gen_burstlen_dest_out(dp_gen_secondary_i_gen_burstlen_dest_out),
    .gen_thread_out(dp_gen_secondary_i_gen_thread_out),
    .gen_mcast_out(dp_gen_secondary_i_gen_mcast_out),
    .gen_data_out(dp_gen_secondary_i_gen_data_out),
    .log_out(dp_gen_secondary_i_log_out),
    .log_valid_out(dp_gen_secondary_i_log_valid_out));
  /* ../../HW/src/dp/dp_fetch.vhd:1256:4  */
  assign n11633_o = n11575_o[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1256:4  */
  assign n11634_o = n11575_o[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1256:4  */
  assign n11635_o = n11575_o[72:48];
  /* ../../HW/src/dp/dp_fetch.vhd:1824:5  */
  assign n11636_o = n11575_o[97:73];
  /* ../../HW/src/dp/dp_fetch.vhd:1824:5  */
  assign n11637_o = n11575_o[121:98];
  /* ../../HW/src/dp/dp_fetch.vhd:1824:5  */
  assign n11638_o = n11575_o[145:122];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11639_o = n11575_o[170:146];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11640_o = n11575_o[195:171];
  /* ../../HW/src/dp/dp_fetch.vhd:1352:5  */
  assign n11641_o = n11575_o[219:196];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11642_o = n11575_o[243:220];
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n11643_o = n11575_o[268:244];
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n11644_o = n11575_o[293:269];
  /* ../../HW/src/dp/dp_fetch.vhd:1862:5  */
  assign n11645_o = n11575_o[317:294];
  /* ../../HW/src/dp/dp_fetch.vhd:1862:5  */
  assign n11646_o = n11575_o[341:318];
  /* ../../HW/src/dp/dp_fetch.vhd:1862:5  */
  assign n11647_o = n11575_o[366:342];
  /* ../../HW/src/dp/dp_fetch.vhd:1352:5  */
  assign n11648_o = n11575_o[391:367];
  /* ../../HW/src/dp/dp_fetch.vhd:1285:5  */
  assign n11649_o = n11575_o[415:392];
  /* ../../HW/src/dp/dp_fetch.vhd:1706:1  */
  assign n11650_o = n11575_o[439:416];
  /* ../../HW/src/dp/dp_fetch.vhd:1706:1  */
  assign n11651_o = n11575_o[464:440];
  /* ../../HW/src/dp/dp_fetch.vhd:1706:1  */
  assign n11652_o = n11575_o[489:465];
  /* ../../HW/src/dp/dp_fetch.vhd:1706:1  */
  assign n11653_o = n11575_o[514:490];
  /* ../../HW/src/dp/dp_fetch.vhd:1807:5  */
  assign n11654_o = n11575_o[539:515];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11655_o = n11575_o[564:540];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11656_o = n11575_o[567:565];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11657_o = n11575_o[592:568];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11658_o = n11575_o[624:593];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11659_o = n11575_o[648:625];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n11660_o = n11575_o[672:649];
  assign n11661_o = n11575_o[673];
  assign n11662_o = n11575_o[675:674];
  assign n11663_o = n11575_o[676];
  assign n11664_o = n11575_o[700:677];
  assign n11665_o = n11575_o[706:701];
  assign n11666_o = n11575_o[722:707];
  assign n11667_o = n11575_o[723];
  assign n11668_o = n11575_o[725:724];
  assign n11669_o = n11575_o[727:726];
  assign n11670_o = n11575_o[751:728];
  assign n11671_o = n11575_o[775:752];
  assign n11672_o = n11576_o[23:0];
  assign n11673_o = n11576_o[47:24];
  assign n11674_o = n11576_o[72:48];
  assign n11675_o = n11576_o[97:73];
  assign n11676_o = n11576_o[121:98];
  assign n11677_o = n11576_o[145:122];
  assign n11678_o = n11576_o[170:146];
  assign n11679_o = n11576_o[195:171];
  assign n11680_o = n11576_o[219:196];
  assign n11681_o = n11576_o[243:220];
  assign n11682_o = n11576_o[268:244];
  assign n11683_o = n11576_o[293:269];
  assign n11684_o = n11576_o[317:294];
  assign n11685_o = n11576_o[341:318];
  assign n11686_o = n11576_o[366:342];
  assign n11687_o = n11576_o[391:367];
  assign n11688_o = n11576_o[415:392];
  assign n11689_o = n11576_o[439:416];
  assign n11690_o = n11576_o[464:440];
  assign n11691_o = n11576_o[489:465];
  assign n11692_o = n11576_o[514:490];
  assign n11693_o = n11576_o[539:515];
  assign n11694_o = n11576_o[564:540];
  assign n11695_o = n11576_o[567:565];
  assign n11696_o = n11576_o[592:568];
  assign n11697_o = n11576_o[624:593];
  assign n11698_o = n11576_o[648:625];
  assign n11699_o = n11576_o[672:649];
  assign n11700_o = n11576_o[673];
  assign n11701_o = n11576_o[675:674];
  assign n11702_o = n11576_o[676];
  assign n11703_o = n11576_o[700:677];
  assign n11704_o = n11576_o[706:701];
  assign n11705_o = n11576_o[722:707];
  assign n11706_o = n11576_o[723];
  assign n11707_o = n11576_o[725:724];
  assign n11708_o = n11576_o[727:726];
  assign n11709_o = n11576_o[751:728];
  assign n11710_o = n11576_o[775:752];
  assign n11711_o = n11580_o[23:0];
  assign n11712_o = n11580_o[47:24];
  assign n11713_o = n11580_o[72:48];
  assign n11714_o = n11580_o[97:73];
  assign n11715_o = n11580_o[121:98];
  assign n11716_o = n11580_o[145:122];
  assign n11717_o = n11580_o[170:146];
  assign n11718_o = n11580_o[195:171];
  assign n11719_o = n11580_o[219:196];
  assign n11720_o = n11580_o[243:220];
  assign n11721_o = n11580_o[268:244];
  assign n11722_o = n11580_o[293:269];
  assign n11723_o = n11580_o[317:294];
  assign n11724_o = n11580_o[341:318];
  assign n11725_o = n11580_o[366:342];
  assign n11726_o = n11580_o[391:367];
  assign n11727_o = n11580_o[415:392];
  assign n11728_o = n11580_o[439:416];
  assign n11729_o = n11580_o[464:440];
  assign n11730_o = n11580_o[489:465];
  assign n11731_o = n11580_o[514:490];
  assign n11732_o = n11580_o[539:515];
  assign n11733_o = n11580_o[564:540];
  assign n11734_o = n11580_o[567:565];
  assign n11735_o = n11580_o[592:568];
  assign n11736_o = n11580_o[624:593];
  assign n11737_o = n11580_o[648:625];
  assign n11738_o = n11580_o[672:649];
  assign n11739_o = n11580_o[673];
  assign n11740_o = n11580_o[675:674];
  assign n11741_o = n11580_o[676];
  assign n11742_o = n11580_o[700:677];
  assign n11743_o = n11580_o[706:701];
  assign n11744_o = n11580_o[722:707];
  assign n11745_o = n11580_o[723];
  assign n11746_o = n11580_o[725:724];
  assign n11747_o = n11580_o[727:726];
  assign n11748_o = n11580_o[751:728];
  assign n11749_o = n11580_o[775:752];
  assign n11750_o = n11581_o[23:0];
  assign n11751_o = n11581_o[47:24];
  assign n11752_o = n11581_o[72:48];
  assign n11753_o = n11581_o[97:73];
  assign n11754_o = n11581_o[121:98];
  assign n11755_o = n11581_o[145:122];
  assign n11756_o = n11581_o[170:146];
  assign n11757_o = n11581_o[195:171];
  assign n11758_o = n11581_o[219:196];
  assign n11759_o = n11581_o[243:220];
  assign n11760_o = n11581_o[268:244];
  assign n11761_o = n11581_o[293:269];
  assign n11762_o = n11581_o[317:294];
  assign n11763_o = n11581_o[341:318];
  assign n11764_o = n11581_o[366:342];
  assign n11765_o = n11581_o[391:367];
  assign n11766_o = n11581_o[415:392];
  assign n11767_o = n11581_o[439:416];
  assign n11768_o = n11581_o[464:440];
  assign n11769_o = n11581_o[489:465];
  assign n11770_o = n11581_o[514:490];
  assign n11771_o = n11581_o[539:515];
  assign n11772_o = n11581_o[564:540];
  assign n11773_o = n11581_o[567:565];
  assign n11774_o = n11581_o[592:568];
  assign n11775_o = n11581_o[624:593];
  assign n11776_o = n11581_o[648:625];
  assign n11777_o = n11581_o[672:649];
  assign n11778_o = n11581_o[673];
  assign n11779_o = n11581_o[675:674];
  assign n11780_o = n11581_o[676];
  assign n11781_o = n11581_o[700:677];
  assign n11782_o = n11581_o[706:701];
  assign n11783_o = n11581_o[722:707];
  assign n11784_o = n11581_o[723];
  assign n11785_o = n11581_o[725:724];
  assign n11786_o = n11581_o[727:726];
  assign n11787_o = n11581_o[751:728];
  assign n11788_o = n11581_o[775:752];
  assign n11856_o = {dp_gen_secondary_i_n11572, dp_gen_primary_i_n11288};
endmodule

module dp_fetch_0_3_3
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [11:0] bus_waddr_in,
   input  [11:0] bus_raddr_in,
   input  bus_write_in,
   input  bus_read_in,
   input  [31:0] bus_writedata_in,
   input  [1:0] ready_in,
   input  [47:0] pcore_sink_counter_in,
   input  [47:0] sram_sink_counter_in,
   input  [23:0] ddr_sink_counter_in,
   input  [1:0] task_busy_in,
   input  task_ready_in,
   input  [31:0] log1_in,
   input  log1_valid_in,
   input  [31:0] log2_in,
   input  log2_valid_in,
   input  [2:0] pcore_read_pending_p0_in,
   input  [2:0] sram_read_pending_p0_in,
   input  [2:0] ddr_read_pending_p0_in,
   input  [2:0] pcore_read_pending_p1_in,
   input  [2:0] sram_read_pending_p1_in,
   input  [2:0] ddr_read_pending_p1_in,
   input  ddr_tx_busy_in,
   output [31:0] bus_readdata_out,
   output bus_readdatavalid_out,
   output bus_writewait_out,
   output bus_readwait_out,
   output [1:0] instruction_valid_out,
   output [2:0] instruction_out_opcode,
   output [3:0] instruction_out_condition,
   output instruction_out_vm,
   output [775:0] instruction_out_source,
   output [1:0] instruction_out_source_bus_id,
   output [1:0] instruction_out_source_data_type,
   output [775:0] instruction_out_dest,
   output [1:0] instruction_out_dest_bus_id,
   output [1:0] instruction_out_dest_data_type,
   output [5:0] instruction_out_mcast,
   output [23:0] instruction_out_count,
   output [15:0] instruction_out_data,
   output instruction_out_repeat,
   output instruction_out_source_addr_mode,
   output instruction_out_dest_addr_mode,
   output instruction_out_stream_process,
   output [1:0] instruction_out_stream_process_id,
   output [2:0] pre_instruction_out_opcode,
   output [3:0] pre_instruction_out_condition,
   output pre_instruction_out_vm,
   output [775:0] pre_instruction_out_source,
   output [1:0] pre_instruction_out_source_bus_id,
   output [1:0] pre_instruction_out_source_data_type,
   output [775:0] pre_instruction_out_dest,
   output [1:0] pre_instruction_out_dest_bus_id,
   output [1:0] pre_instruction_out_dest_data_type,
   output [5:0] pre_instruction_out_mcast,
   output [23:0] pre_instruction_out_count,
   output [15:0] pre_instruction_out_data,
   output pre_instruction_out_repeat,
   output pre_instruction_out_source_addr_mode,
   output pre_instruction_out_dest_addr_mode,
   output pre_instruction_out_stream_process,
   output [1:0] pre_instruction_out_stream_process_id,
   output [10:0] task_start_addr_out,
   output task_pending_out,
   output task_out,
   output task_vm_out,
   output [4:0] task_pcore_out,
   output task_lockstep_out,
   output [3:0] task_tid_mask_out,
   output [27:0] task_iregister_auto_out,
   output [1:0] task_data_model_out,
   output indication_avail_out);
  wire [2:0] n7776_o;
  wire [3:0] n7777_o;
  wire n7778_o;
  wire [775:0] n7779_o;
  wire [1:0] n7780_o;
  wire [1:0] n7781_o;
  wire [775:0] n7782_o;
  wire [1:0] n7783_o;
  wire [1:0] n7784_o;
  wire [5:0] n7785_o;
  wire [23:0] n7786_o;
  wire [15:0] n7787_o;
  wire n7788_o;
  wire n7789_o;
  wire n7790_o;
  wire n7791_o;
  wire [1:0] n7792_o;
  wire [2:0] n7794_o;
  wire [3:0] n7795_o;
  wire n7796_o;
  wire [775:0] n7797_o;
  wire [1:0] n7798_o;
  wire [1:0] n7799_o;
  wire [775:0] n7800_o;
  wire [1:0] n7801_o;
  wire [1:0] n7802_o;
  wire [5:0] n7803_o;
  wire [23:0] n7804_o;
  wire [15:0] n7805_o;
  wire n7806_o;
  wire n7807_o;
  wire n7808_o;
  wire n7809_o;
  wire [1:0] n7810_o;
  wire [7:0] fifo_avail;
  wire match;
  wire [1619:0] irec;
  wire [96:0] irec_generic;
  wire [1619:0] orec;
  wire [3239:0] orecs;
  wire [96:0] orec_generic;
  wire [1517:0] data;
  wire [1517:0] q1;
  wire [1517:0] q2;
  wire rdreq;
  wire [1:0] rdreqs;
  wire wreq;
  wire wreq_all;
  wire full;
  wire ready;
  wire ready_which;
  wire [1:0] ready2;
  wire valid;
  wire [1:0] valids;
  wire [4:0] wregno;
  wire [4:0] rregno;
  wire [47:0] pcore_sink_counter_r;
  wire [47:0] sram_sink_counter_r;
  wire [23:0] ddr_sink_counter_r;
  wire [1:0] sink_pcore_busy_r;
  wire [1:0] sink_sram_busy_r;
  wire sink_ddr_busy_r;
  wire [1:0] pcore_source_busy_r;
  wire [1:0] sram_source_busy_r;
  wire ddr_source_busy_r;
  wire log_enable_r;
  wire print_indication_r;
  wire print_indication_rr;
  wire [63:0] print_param_r;
  wire [63:0] print_param_rr;
  wire wreq2;
  wire wreq2_indication;
  wire [2:0] pcore_read_pending;
  wire [2:0] sram_read_pending;
  wire [2:0] ddr_read_pending;
  wire indication_full_r;
  wire indication_rdreq;
  wire [66:0] in_indication;
  wire [66:0] indication;
  wire [7:0] indication_rdusedw;
  wire [7:0] indication_wrusedw;
  wire [63:0] indication_parm_r;
  wire [31:0] indication_r;
  wire indication_sync_r;
  wire [31:0] bus_readdata_r;
  wire [1:0] instruction_valid_r;
  wire [1:0] instruction_valid_rr;
  wire [1619:0] instruction_r;
  wire [1619:0] instruction_rr;
  wire [1619:0] instruction;
  wire [63:0] log_status_last_r;
  wire [63:0] log_write;
  wire [63:0] log_read;
  wire [31:0] log_readtime_r;
  wire log_rdreq;
  wire log_empty;
  wire log_full;
  wire [31:0] log_time_r;
  wire log_wrreq;
  wire log_wrreq2;
  wire load;
  wire load_r;
  wire [3:0] load_busid_r;
  wire [3:0] dp_var_waddress;
  wire [3:0] dp_var_raddress;
  wire [775:0] dp_var_write;
  wire [775:0] dp_var_read;
  wire dp_var_we;
  wire [775:0] dp_var_template;
  wire task2;
  wire waitrequest;
  wire [3:0] source_bus_id_r;
  wire [1:0] source_vm_r;
  wire [3:0] dest_bus_id_r;
  wire outoforderok;
  wire [15:0] new_cmd_is_safe_r;
  wire [3:0] condition_vm0_busy_r;
  wire [3:0] condition_vm1_busy_r;
  wire curr_vm_r;
  wire [1:0] pcore_sink_busy_r;
  wire [1:0] sram_sink_busy_r;
  wire ddr_sink_busy_r;
  wire [5:0] wregno2;
  wire [5:0] wregno2_r;
  reg [775:0] src_template_r;
  reg [775:0] dest_template_r;
  reg [775:0] template_r;
  wire pause;
  wire [1:0] pauses;
  wire [10:0] task_start_addr;
  wire [4:0] task_pcore;
  wire [3:0] task_tid_mask;
  wire [1:0] task_data_model;
  wire [27:0] task_iregister_auto;
  wire task_lockstep;
  wire \task ;
  wire task_vm;
  wire [10:0] task_start_addr_r;
  reg [4:0] task_pcore_r;
  reg [3:0] task_tid_mask_r;
  wire [1:0] task_data_model_r;
  wire [27:0] task_iregister_auto_r;
  wire task_lockstep_r;
  wire task_r;
  wire task_vm_r;
  wire [11:0] bus_waddr_r;
  wire [11:0] bus_raddr_r;
  wire bus_write_r;
  wire bus_read_r;
  wire [31:0] bus_writedata_r;
  wire rden_r;
  wire [1:0] avail;
  wire indication_empty;
  wire n7826_o;
  wire n7827_o;
  wire n7828_o;
  wire n7829_o;
  wire n7830_o;
  wire n7831_o;
  wire n7832_o;
  wire n7833_o;
  wire n7834_o;
  wire n7835_o;
  wire n7836_o;
  wire n7837_o;
  wire n7838_o;
  wire n7839_o;
  wire n7840_o;
  wire n7841_o;
  wire n7842_o;
  wire [1:0] n7843_o;
  wire [1:0] n7844_o;
  wire [1:0] n7845_o;
  wire [1:0] n7846_o;
  wire n7848_o;
  wire n7849_o;
  wire [4:0] n7850_o;
  wire n7852_o;
  wire n7853_o;
  wire n7854_o;
  wire n7855_o;
  localparam n7857_o = 1'b0;
  wire n7860_o;
  wire n7861_o;
  wire n7863_o;
  wire n7864_o;
  wire n7865_o;
  wire [31:0] n7869_o;
  wire [29:0] n7871_o;
  wire n7872_o;
  wire n7873_o;
  wire n7874_o;
  wire n7875_o;
  wire n7876_o;
  wire n7877_o;
  wire n7878_o;
  wire n7879_o;
  wire n7880_o;
  wire n7881_o;
  wire [19:0] n7882_o;
  localparam [31:0] n7883_o = 32'b00000000000000000000000000000000;
  wire [29:0] n7885_o;
  wire [11:0] n7886_o;
  wire [11:0] n7887_o;
  wire n7888_o;
  wire n7891_o;
  wire [31:0] n7892_o;
  wire [31:0] n7893_o;
  wire n7895_o;
  wire [31:0] n7896_o;
  wire n7898_o;
  wire [63:0] n7899_o;
  wire [63:0] n7900_o;
  wire [63:0] n7901_o;
  wire n7903_o;
  wire n7905_o;
  wire n7906_o;
  wire n7907_o;
  wire [63:0] log_fifo_i_n7908;
  wire log_fifo_i_n7911;
  wire log_fifo_i_n7912;
  wire [63:0] log_fifo_i_q_out;
  wire [7:0] log_fifo_i_ravail_out;
  wire [7:0] log_fifo_i_wused_out;
  wire log_fifo_i_empty_out;
  wire log_fifo_i_full_out;
  wire log_fifo_i_almost_full_out;
  wire n7924_o;
  wire n7925_o;
  wire n7926_o;
  wire n7927_o;
  wire [1517:0] fifo_i_n7929;
  wire [1517:0] fifo_i_n7930;
  wire n7931_o;
  wire n7932_o;
  wire fifo_i_n7933;
  wire fifo_i_n7934;
  wire fifo_i_n7935;
  wire [7:0] fifo_i_n7936;
  wire [1517:0] fifo_i_readdata1_out;
  wire [1517:0] fifo_i_readdata2_out;
  wire fifo_i_valid1_out;
  wire fifo_i_valid2_out;
  wire fifo_i_full_out;
  wire [7:0] fifo_i_fifo_avail_out;
  wire [775:0] gen1_ram_i_n7949;
  wire [775:0] gen1_ram_i_q_b;
  wire [23:0] n7959_o;
  wire [23:0] n7962_o;
  wire [24:0] n7964_o;
  wire [24:0] n7966_o;
  wire [23:0] n7968_o;
  wire [23:0] n7970_o;
  wire [24:0] n7972_o;
  wire [24:0] n7974_o;
  wire [23:0] n7976_o;
  wire [23:0] n7978_o;
  wire [24:0] n7980_o;
  wire [24:0] n7982_o;
  wire [23:0] n7984_o;
  wire [23:0] n7986_o;
  wire [24:0] n7988_o;
  wire [24:0] n7990_o;
  wire [23:0] n7992_o;
  wire [23:0] n7994_o;
  wire [24:0] n7996_o;
  wire [24:0] n7998_o;
  wire [24:0] n8000_o;
  wire [24:0] n8002_o;
  wire [24:0] n8004_o;
  wire [2:0] n8006_o;
  wire [24:0] n8008_o;
  wire [31:0] n8010_o;
  wire [23:0] n8012_o;
  wire [23:0] n8014_o;
  wire n8016_o;
  wire [1:0] n8018_o;
  wire n8020_o;
  wire [23:0] n8022_o;
  wire [5:0] n8024_o;
  wire [15:0] n8026_o;
  wire n8028_o;
  wire [1:0] n8030_o;
  wire [1:0] n8032_o;
  wire [23:0] n8034_o;
  wire [23:0] n8036_o;
  wire [775:0] n8037_o;
  wire [23:0] n8045_o;
  wire [23:0] n8048_o;
  wire [24:0] n8050_o;
  wire [24:0] n8052_o;
  wire [23:0] n8054_o;
  wire [23:0] n8056_o;
  wire [24:0] n8058_o;
  wire [24:0] n8060_o;
  wire [23:0] n8062_o;
  wire [23:0] n8064_o;
  wire [24:0] n8066_o;
  wire [24:0] n8068_o;
  wire [23:0] n8070_o;
  wire [23:0] n8072_o;
  wire [24:0] n8074_o;
  wire [24:0] n8076_o;
  wire [23:0] n8078_o;
  wire [23:0] n8080_o;
  wire [24:0] n8082_o;
  wire [24:0] n8084_o;
  wire [24:0] n8086_o;
  wire [24:0] n8088_o;
  wire [24:0] n8090_o;
  wire [2:0] n8092_o;
  wire [24:0] n8094_o;
  wire [31:0] n8096_o;
  wire [23:0] n8098_o;
  wire [23:0] n8100_o;
  wire n8102_o;
  wire [1:0] n8104_o;
  wire n8106_o;
  wire [23:0] n8108_o;
  wire [5:0] n8110_o;
  wire [15:0] n8112_o;
  wire n8114_o;
  wire [1:0] n8116_o;
  wire [1:0] n8118_o;
  wire [23:0] n8120_o;
  wire [23:0] n8122_o;
  wire [775:0] n8123_o;
  wire [3:0] n8124_o;
  wire n8125_o;
  wire [3:0] n8126_o;
  wire [2:0] n8127_o;
  wire [3:0] n8128_o;
  wire [2:0] n8129_o;
  wire [63:0] n8130_o;
  wire [66:0] n8131_o;
  wire [66:0] indication_i_n8132;
  wire [7:0] indication_i_n8133;
  wire [7:0] indication_i_n8134;
  wire indication_i_n8135;
  wire [66:0] indication_i_q_out;
  wire [7:0] indication_i_ravail_out;
  wire [7:0] indication_i_wused_out;
  wire indication_i_empty_out;
  wire indication_i_full_out;
  wire indication_i_almost_full_out;
  wire [2:0] n8149_o;
  wire [2:0] n8150_o;
  wire [2:0] n8151_o;
  wire [4:0] n8152_o;
  wire [5:0] n8153_o;
  wire [5:0] n8154_o;
  wire [4:0] n8155_o;
  wire [2:0] n8166_o;
  wire [3:0] n8169_o;
  wire n8171_o;
  wire [775:0] n8173_o;
  wire [23:0] n8174_o;
  wire [775:0] n8176_o;
  wire [23:0] n8177_o;
  wire [775:0] n8179_o;
  wire [24:0] n8180_o;
  wire [775:0] n8182_o;
  wire [24:0] n8183_o;
  wire [775:0] n8185_o;
  wire [23:0] n8186_o;
  wire [775:0] n8188_o;
  wire [23:0] n8189_o;
  wire [775:0] n8191_o;
  wire [24:0] n8192_o;
  wire [775:0] n8194_o;
  wire [24:0] n8195_o;
  wire [775:0] n8197_o;
  wire [23:0] n8198_o;
  wire [775:0] n8200_o;
  wire [23:0] n8201_o;
  wire [775:0] n8203_o;
  wire [24:0] n8204_o;
  wire [775:0] n8206_o;
  wire [24:0] n8207_o;
  wire [775:0] n8209_o;
  wire [23:0] n8210_o;
  wire [775:0] n8212_o;
  wire [23:0] n8213_o;
  wire [775:0] n8215_o;
  wire [24:0] n8216_o;
  wire [775:0] n8218_o;
  wire [24:0] n8219_o;
  wire [775:0] n8221_o;
  wire [23:0] n8222_o;
  wire [775:0] n8224_o;
  wire [23:0] n8225_o;
  wire [775:0] n8227_o;
  wire [24:0] n8228_o;
  wire [775:0] n8230_o;
  wire [24:0] n8231_o;
  wire [775:0] n8233_o;
  wire [24:0] n8234_o;
  wire [775:0] n8236_o;
  wire [24:0] n8237_o;
  wire [775:0] n8239_o;
  wire [24:0] n8240_o;
  wire [775:0] n8242_o;
  wire [2:0] n8243_o;
  wire [775:0] n8245_o;
  wire [24:0] n8246_o;
  wire [775:0] n8248_o;
  wire n8249_o;
  wire [775:0] n8251_o;
  wire [1:0] n8252_o;
  wire [775:0] n8254_o;
  wire n8255_o;
  wire [775:0] n8257_o;
  wire [31:0] n8258_o;
  wire [775:0] n8260_o;
  wire [23:0] n8261_o;
  wire [775:0] n8263_o;
  wire [23:0] n8264_o;
  wire [775:0] n8266_o;
  wire [23:0] n8267_o;
  wire [775:0] n8269_o;
  wire [23:0] n8270_o;
  wire [1:0] n8272_o;
  wire [1:0] n8274_o;
  wire [775:0] n8276_o;
  wire [23:0] n8277_o;
  wire [775:0] n8279_o;
  wire [23:0] n8280_o;
  wire [775:0] n8282_o;
  wire [24:0] n8283_o;
  wire [775:0] n8285_o;
  wire [24:0] n8286_o;
  wire [775:0] n8288_o;
  wire [23:0] n8289_o;
  wire [775:0] n8291_o;
  wire [23:0] n8292_o;
  wire [775:0] n8294_o;
  wire [24:0] n8295_o;
  wire [775:0] n8297_o;
  wire [24:0] n8298_o;
  wire [775:0] n8300_o;
  wire [23:0] n8301_o;
  wire [775:0] n8303_o;
  wire [23:0] n8304_o;
  wire [775:0] n8306_o;
  wire [24:0] n8307_o;
  wire [775:0] n8309_o;
  wire [24:0] n8310_o;
  wire [775:0] n8312_o;
  wire [23:0] n8313_o;
  wire [775:0] n8315_o;
  wire [23:0] n8316_o;
  wire [775:0] n8318_o;
  wire [24:0] n8319_o;
  wire [775:0] n8321_o;
  wire [24:0] n8322_o;
  wire [775:0] n8324_o;
  wire [23:0] n8325_o;
  wire [775:0] n8327_o;
  wire [23:0] n8328_o;
  wire [775:0] n8330_o;
  wire [24:0] n8331_o;
  wire [775:0] n8333_o;
  wire [24:0] n8334_o;
  wire [775:0] n8336_o;
  wire [24:0] n8337_o;
  wire [775:0] n8339_o;
  wire [24:0] n8340_o;
  wire [775:0] n8342_o;
  wire [24:0] n8343_o;
  wire [775:0] n8345_o;
  wire [2:0] n8346_o;
  wire [775:0] n8348_o;
  wire [24:0] n8349_o;
  wire [775:0] n8351_o;
  wire n8352_o;
  wire [775:0] n8354_o;
  wire [1:0] n8355_o;
  wire [775:0] n8357_o;
  wire n8358_o;
  wire [775:0] n8360_o;
  wire [31:0] n8361_o;
  wire [775:0] n8363_o;
  wire [23:0] n8364_o;
  wire [775:0] n8366_o;
  wire [23:0] n8367_o;
  wire [775:0] n8369_o;
  wire [23:0] n8370_o;
  wire [775:0] n8372_o;
  wire [23:0] n8373_o;
  wire [1:0] n8375_o;
  wire [1:0] n8377_o;
  wire [5:0] n8379_o;
  wire [23:0] n8381_o;
  wire [15:0] n8383_o;
  wire n8385_o;
  wire n8387_o;
  wire n8389_o;
  wire n8391_o;
  wire [1:0] n8393_o;
  wire [1517:0] n8394_o;
  wire [2:0] n8395_o;
  wire n8397_o;
  wire [1517:0] n8398_o;
  wire [2:0] n8406_o;
  wire [3:0] n8407_o;
  wire [6:0] n8408_o;
  wire n8409_o;
  wire [7:0] n8410_o;
  wire [24:0] n8411_o;
  wire [32:0] n8412_o;
  wire [63:0] n8413_o;
  wire [96:0] n8414_o;
  wire [1517:0] n8416_o;
  wire [2:0] n8425_o;
  localparam [1619:0] n8426_o = 1620'bX;
  wire [3:0] n8428_o;
  wire n8430_o;
  wire [23:0] n8432_o;
  wire [23:0] n8434_o;
  wire [24:0] n8436_o;
  wire [24:0] n8438_o;
  wire [23:0] n8440_o;
  wire [23:0] n8442_o;
  wire [24:0] n8444_o;
  wire [24:0] n8446_o;
  wire [23:0] n8448_o;
  wire [23:0] n8450_o;
  wire [24:0] n8452_o;
  wire [24:0] n8454_o;
  wire [23:0] n8456_o;
  wire [23:0] n8458_o;
  wire [24:0] n8460_o;
  wire [24:0] n8462_o;
  wire [23:0] n8464_o;
  wire [23:0] n8466_o;
  wire [24:0] n8468_o;
  wire [24:0] n8470_o;
  wire [24:0] n8472_o;
  wire [24:0] n8474_o;
  wire [24:0] n8476_o;
  wire [2:0] n8478_o;
  wire [24:0] n8480_o;
  wire n8482_o;
  wire [1:0] n8485_o;
  wire n8487_o;
  wire [31:0] n8489_o;
  wire [23:0] n8491_o;
  wire [23:0] n8493_o;
  wire [23:0] n8494_o;
  wire [50:0] n8496_o;
  wire [23:0] n8497_o;
  wire [1:0] n8499_o;
  wire [1:0] n8501_o;
  wire [23:0] n8503_o;
  wire [23:0] n8505_o;
  wire [24:0] n8507_o;
  wire [24:0] n8509_o;
  wire [23:0] n8511_o;
  wire [23:0] n8513_o;
  wire [24:0] n8515_o;
  wire [24:0] n8517_o;
  wire [23:0] n8519_o;
  wire [23:0] n8521_o;
  wire [24:0] n8523_o;
  wire [24:0] n8525_o;
  wire [23:0] n8527_o;
  wire [23:0] n8529_o;
  wire [24:0] n8531_o;
  wire [24:0] n8533_o;
  wire [23:0] n8535_o;
  wire [23:0] n8537_o;
  wire [24:0] n8539_o;
  wire [24:0] n8541_o;
  wire [24:0] n8543_o;
  wire [24:0] n8545_o;
  wire [24:0] n8547_o;
  wire [2:0] n8549_o;
  wire [24:0] n8551_o;
  wire n8553_o;
  wire [1:0] n8556_o;
  wire n8558_o;
  wire [31:0] n8560_o;
  wire [23:0] n8562_o;
  wire [23:0] n8564_o;
  wire [23:0] n8565_o;
  wire [50:0] n8567_o;
  wire [23:0] n8568_o;
  wire [1:0] n8570_o;
  wire [1:0] n8572_o;
  wire [5:0] n8574_o;
  wire [23:0] n8576_o;
  wire [15:0] n8578_o;
  wire n8580_o;
  wire n8582_o;
  wire n8584_o;
  wire n8586_o;
  wire [1:0] n8588_o;
  wire [1619:0] n8589_o;
  wire [2:0] n8597_o;
  localparam [1619:0] n8598_o = 1620'bX;
  wire [3:0] n8600_o;
  wire n8602_o;
  wire [23:0] n8604_o;
  wire [23:0] n8606_o;
  wire [24:0] n8608_o;
  wire [24:0] n8610_o;
  wire [23:0] n8612_o;
  wire [23:0] n8614_o;
  wire [24:0] n8616_o;
  wire [24:0] n8618_o;
  wire [23:0] n8620_o;
  wire [23:0] n8622_o;
  wire [24:0] n8624_o;
  wire [24:0] n8626_o;
  wire [23:0] n8628_o;
  wire [23:0] n8630_o;
  wire [24:0] n8632_o;
  wire [24:0] n8634_o;
  wire [23:0] n8636_o;
  wire [23:0] n8638_o;
  wire [24:0] n8640_o;
  wire [24:0] n8642_o;
  wire [24:0] n8644_o;
  wire [24:0] n8646_o;
  wire [24:0] n8648_o;
  wire [2:0] n8650_o;
  wire [24:0] n8652_o;
  wire n8654_o;
  wire [1:0] n8657_o;
  wire n8659_o;
  wire [31:0] n8661_o;
  wire [23:0] n8663_o;
  wire [23:0] n8665_o;
  wire [23:0] n8666_o;
  wire [50:0] n8668_o;
  wire [23:0] n8669_o;
  wire [1:0] n8671_o;
  wire [1:0] n8673_o;
  wire [23:0] n8675_o;
  wire [23:0] n8677_o;
  wire [24:0] n8679_o;
  wire [24:0] n8681_o;
  wire [23:0] n8683_o;
  wire [23:0] n8685_o;
  wire [24:0] n8687_o;
  wire [24:0] n8689_o;
  wire [23:0] n8691_o;
  wire [23:0] n8693_o;
  wire [24:0] n8695_o;
  wire [24:0] n8697_o;
  wire [23:0] n8699_o;
  wire [23:0] n8701_o;
  wire [24:0] n8703_o;
  wire [24:0] n8705_o;
  wire [23:0] n8707_o;
  wire [23:0] n8709_o;
  wire [24:0] n8711_o;
  wire [24:0] n8713_o;
  wire [24:0] n8715_o;
  wire [24:0] n8717_o;
  wire [24:0] n8719_o;
  wire [2:0] n8721_o;
  wire [24:0] n8723_o;
  wire n8725_o;
  wire [1:0] n8728_o;
  wire n8730_o;
  wire [31:0] n8732_o;
  wire [23:0] n8734_o;
  wire [23:0] n8736_o;
  wire [23:0] n8737_o;
  wire [50:0] n8739_o;
  wire [23:0] n8740_o;
  wire [1:0] n8742_o;
  wire [1:0] n8744_o;
  wire [5:0] n8746_o;
  wire [23:0] n8748_o;
  wire [15:0] n8750_o;
  wire n8752_o;
  wire n8754_o;
  wire n8756_o;
  wire n8758_o;
  wire [1:0] n8760_o;
  wire [1619:0] n8761_o;
  wire [2:0] n8769_o;
  wire [3:0] n8772_o;
  wire n8774_o;
  wire [24:0] n8776_o;
  wire [63:0] n8778_o;
  wire [96:0] n8779_o;
  wire [1:0] n8781_o;
  wire [1:0] n8782_o;
  wire [1:0] n8783_o;
  wire [5:0] n8784_o;
  wire [23:0] n8785_o;
  wire [15:0] n8786_o;
  wire n8787_o;
  wire [2:0] n8795_o;
  wire [3:0] n8798_o;
  wire n8808_o;
  wire n8811_o;
  wire n8813_o;
  wire [1:0] n8815_o;
  wire [1619:0] n8819_o;
  wire [2:0] n8827_o;
  wire [3:0] n8830_o;
  wire [24:0] n8833_o;
  wire [96:0] n8835_o;
  wire n8838_o;
  wire n8839_o;
  wire n8840_o;
  wire n8842_o;
  wire n8844_o;
  wire n8845_o;
  wire [2:0] n8846_o;
  wire n8848_o;
  wire n8849_o;
  wire n8850_o;
  wire n8853_o;
  wire n8854_o;
  wire [2:0] n8855_o;
  wire n8857_o;
  wire n8858_o;
  wire n8859_o;
  wire [2:0] n8863_o;
  wire n8865_o;
  wire n8866_o;
  wire n8867_o;
  wire [1:0] n8868_o;
  wire [1:0] n8869_o;
  wire n8870_o;
  wire [1:0] n8871_o;
  wire [1:0] n8872_o;
  wire n8873_o;
  wire n8874_o;
  wire n8875_o;
  wire n8876_o;
  wire n8877_o;
  wire n8878_o;
  wire n8879_o;
  wire [1:0] n8880_o;
  wire [1:0] n8881_o;
  wire n8882_o;
  wire [1:0] n8883_o;
  wire [1:0] n8884_o;
  wire n8885_o;
  wire n8886_o;
  wire n8887_o;
  wire n8888_o;
  wire n8889_o;
  wire n8890_o;
  wire n8892_o;
  wire n8895_o;
  wire n8896_o;
  wire n8898_o;
  wire n8900_o;
  wire n8902_o;
  wire n8906_o;
  wire n8907_o;
  wire n8908_o;
  wire n8909_o;
  wire n8913_o;
  wire n8914_o;
  wire n8915_o;
  wire n8916_o;
  wire n8917_o;
  wire n8918_o;
  wire n8922_o;
  wire n8924_o;
  wire n8926_o;
  wire n8947_o;
  wire [31:0] n8950_o;
  wire n8951_o;
  wire n8953_o;
  wire [31:0] n8954_o;
  wire n8956_o;
  wire n8959_o;
  wire n8961_o;
  wire [31:0] n8962_o;
  wire n8964_o;
  wire n8967_o;
  wire n8968_o;
  wire [31:0] n8969_o;
  wire [31:0] n8971_o;
  wire [31:0] n8972_o;
  wire n8974_o;
  wire [31:0] n8976_o;
  wire n8979_o;
  wire [31:0] n8980_o;
  wire [31:0] n8981_o;
  wire n8983_o;
  wire [31:0] n8984_o;
  wire [31:0] n8985_o;
  wire [31:0] n8986_o;
  wire n8988_o;
  wire [31:0] n8989_o;
  wire [31:0] n8990_o;
  wire n8992_o;
  wire [31:0] n8993_o;
  wire [31:0] n8994_o;
  wire n8996_o;
  wire [31:0] n8997_o;
  wire [31:0] n8998_o;
  wire [31:0] n8999_o;
  wire n9001_o;
  wire [31:0] n9005_o;
  wire [31:0] n9006_o;
  wire n9008_o;
  wire n9009_o;
  wire n9010_o;
  wire n9014_o;
  wire n9046_o;
  wire n9049_o;
  wire n9051_o;
  wire [775:0] n9052_o;
  wire [775:0] n9054_o;
  wire n9055_o;
  localparam [775:0] n9057_o = 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [775:0] n9058_o;
  wire n9060_o;
  wire n9062_o;
  wire [23:0] n9063_o;
  wire [23:0] n9064_o;
  wire [23:0] n9065_o;
  wire [23:0] n9066_o;
  wire [23:0] n9067_o;
  wire n9069_o;
  wire [23:0] n9070_o;
  wire [23:0] n9071_o;
  wire [23:0] n9072_o;
  wire [23:0] n9073_o;
  wire [23:0] n9074_o;
  wire n9076_o;
  wire [24:0] n9077_o;
  wire [24:0] n9078_o;
  wire [24:0] n9079_o;
  wire [24:0] n9080_o;
  wire [24:0] n9081_o;
  wire n9083_o;
  wire [23:0] n9084_o;
  wire [23:0] n9085_o;
  wire [23:0] n9086_o;
  wire [23:0] n9087_o;
  wire [23:0] n9088_o;
  wire n9090_o;
  wire [23:0] n9091_o;
  wire [23:0] n9092_o;
  wire [23:0] n9093_o;
  wire [23:0] n9094_o;
  wire [23:0] n9095_o;
  wire n9097_o;
  wire [24:0] n9098_o;
  wire [24:0] n9099_o;
  wire [24:0] n9100_o;
  wire [24:0] n9101_o;
  wire [24:0] n9102_o;
  wire n9104_o;
  wire [23:0] n9105_o;
  wire [23:0] n9106_o;
  wire [23:0] n9107_o;
  wire [23:0] n9108_o;
  wire [23:0] n9109_o;
  wire n9111_o;
  wire [23:0] n9112_o;
  wire [23:0] n9113_o;
  wire [23:0] n9114_o;
  wire [23:0] n9115_o;
  wire [23:0] n9116_o;
  wire n9118_o;
  wire [24:0] n9119_o;
  wire [24:0] n9120_o;
  wire [24:0] n9121_o;
  wire [24:0] n9122_o;
  wire [24:0] n9123_o;
  wire n9125_o;
  wire [23:0] n9126_o;
  wire [23:0] n9127_o;
  wire [23:0] n9128_o;
  wire [23:0] n9129_o;
  wire [23:0] n9130_o;
  wire n9132_o;
  wire [23:0] n9133_o;
  wire [23:0] n9134_o;
  wire [23:0] n9135_o;
  wire [23:0] n9136_o;
  wire [23:0] n9137_o;
  wire n9139_o;
  wire [24:0] n9140_o;
  wire [24:0] n9141_o;
  wire [24:0] n9142_o;
  wire [24:0] n9143_o;
  wire [24:0] n9144_o;
  wire n9146_o;
  wire [23:0] n9147_o;
  wire [23:0] n9148_o;
  wire [23:0] n9149_o;
  wire [23:0] n9150_o;
  wire [23:0] n9151_o;
  wire n9153_o;
  wire [23:0] n9154_o;
  wire [23:0] n9155_o;
  wire [23:0] n9156_o;
  wire [23:0] n9157_o;
  wire [23:0] n9158_o;
  wire n9160_o;
  wire [24:0] n9161_o;
  wire [24:0] n9162_o;
  wire [24:0] n9163_o;
  wire [24:0] n9164_o;
  wire [24:0] n9165_o;
  wire n9167_o;
  wire [24:0] n9168_o;
  wire [24:0] n9169_o;
  wire [24:0] n9170_o;
  wire [74:0] n9171_o;
  wire n9177_o;
  wire [24:0] n9178_o;
  wire [24:0] n9179_o;
  wire [24:0] n9180_o;
  wire [24:0] n9181_o;
  wire [24:0] n9182_o;
  wire [24:0] n9183_o;
  wire [24:0] n9184_o;
  wire [24:0] n9185_o;
  wire [24:0] n9186_o;
  wire [24:0] n9187_o;
  wire [24:0] n9188_o;
  wire [24:0] n9189_o;
  wire [24:0] n9190_o;
  wire [24:0] n9191_o;
  wire [24:0] n9192_o;
  wire [24:0] n9193_o;
  wire [24:0] n9194_o;
  wire n9196_o;
  wire [24:0] n9197_o;
  wire [24:0] n9198_o;
  wire n9200_o;
  wire [2:0] n9201_o;
  wire [2:0] n9202_o;
  wire [2:0] n9203_o;
  wire [2:0] n9204_o;
  wire [2:0] n9205_o;
  wire n9207_o;
  wire [31:0] n9208_o;
  wire [31:0] n9209_o;
  wire n9216_o;
  wire [23:0] n9217_o;
  wire [23:0] n9218_o;
  wire [23:0] n9219_o;
  wire [23:0] n9220_o;
  wire [23:0] n9221_o;
  wire n9223_o;
  wire [23:0] n9224_o;
  wire [23:0] n9225_o;
  wire [23:0] n9226_o;
  wire [23:0] n9227_o;
  wire [23:0] n9228_o;
  wire n9230_o;
  wire [23:0] n9231_o;
  wire [23:0] n9232_o;
  wire [23:0] n9233_o;
  wire [23:0] n9234_o;
  wire [23:0] n9235_o;
  wire n9237_o;
  wire [23:0] n9238_o;
  wire [23:0] n9239_o;
  wire [23:0] n9240_o;
  wire [23:0] n9241_o;
  wire [23:0] n9242_o;
  wire n9244_o;
  wire n9245_o;
  wire n9246_o;
  wire [1:0] n9247_o;
  wire [1:0] n9248_o;
  wire n9249_o;
  wire [1:0] n9250_o;
  wire n9252_o;
  wire n9254_o;
  wire n9255_o;
  wire n9256_o;
  wire n9257_o;
  wire n9258_o;
  wire n9259_o;
  wire n9260_o;
  wire n9261_o;
  wire n9262_o;
  wire n9263_o;
  wire n9264_o;
  wire n9265_o;
  wire n9266_o;
  wire n9267_o;
  wire n9268_o;
  wire n9269_o;
  wire n9270_o;
  wire n9271_o;
  wire n9272_o;
  wire n9273_o;
  wire n9274_o;
  wire n9275_o;
  wire n9276_o;
  wire n9277_o;
  wire n9278_o;
  wire n9279_o;
  wire [5:0] n9280_o;
  wire [3:0] n9281_o;
  wire [4:0] n9282_o;
  wire n9283_o;
  wire n9284_o;
  wire n9285_o;
  wire n9286_o;
  wire n9287_o;
  wire n9288_o;
  wire n9289_o;
  wire n9290_o;
  wire n9291_o;
  wire n9292_o;
  wire n9293_o;
  wire n9294_o;
  wire n9295_o;
  wire n9296_o;
  wire n9297_o;
  wire n9298_o;
  wire [3:0] n9299_o;
  wire [3:0] n9300_o;
  wire [3:0] n9301_o;
  wire [3:0] n9302_o;
  wire [5:0] n9303_o;
  wire [5:0] n9304_o;
  wire [5:0] n9305_o;
  wire [5:0] n9306_o;
  wire [4:0] n9307_o;
  wire [4:0] n9308_o;
  wire [4:0] n9309_o;
  wire [4:0] n9310_o;
  wire n9314_o;
  wire [3:0] n9315_o;
  wire [2:0] n9316_o;
  wire [3:0] n9317_o;
  wire [3:0] n9318_o;
  wire n9320_o;
  wire n9321_o;
  wire n9322_o;
  wire n9323_o;
  wire n9324_o;
  wire n9325_o;
  wire n9326_o;
  wire n9327_o;
  wire n9328_o;
  wire n9329_o;
  wire n9330_o;
  wire n9331_o;
  wire n9332_o;
  wire n9333_o;
  wire n9334_o;
  wire n9335_o;
  wire [3:0] n9336_o;
  wire [3:0] n9337_o;
  wire [3:0] n9338_o;
  wire [3:0] n9339_o;
  wire [5:0] n9340_o;
  wire [5:0] n9341_o;
  wire [5:0] n9342_o;
  wire [5:0] n9343_o;
  wire [4:0] n9344_o;
  wire [4:0] n9345_o;
  wire [4:0] n9346_o;
  wire [4:0] n9347_o;
  wire [13:0] n9355_o;
  wire [13:0] n9356_o;
  wire [13:0] n9357_o;
  wire [13:0] n9358_o;
  wire [13:0] n9359_o;
  wire [13:0] n9360_o;
  wire [13:0] n9361_o;
  wire [9:0] n9362_o;
  wire [9:0] n9363_o;
  wire [9:0] n9364_o;
  wire [9:0] n9365_o;
  wire [9:0] n9366_o;
  wire [9:0] n9367_o;
  wire [9:0] n9368_o;
  wire [5:0] n9369_o;
  wire [5:0] n9370_o;
  wire [5:0] n9371_o;
  wire [5:0] n9372_o;
  wire [5:0] n9373_o;
  wire [5:0] n9374_o;
  wire [5:0] n9375_o;
  wire n9379_o;
  wire [24:0] n9380_o;
  wire [24:0] n9381_o;
  wire [24:0] n9382_o;
  wire [24:0] n9383_o;
  wire [24:0] n9384_o;
  wire n9386_o;
  wire [24:0] n9387_o;
  wire [24:0] n9388_o;
  wire [24:0] n9389_o;
  wire [24:0] n9390_o;
  wire [24:0] n9391_o;
  wire n9393_o;
  wire [24:0] n9394_o;
  wire [24:0] n9395_o;
  wire [24:0] n9396_o;
  wire [24:0] n9397_o;
  wire [24:0] n9398_o;
  wire n9400_o;
  wire [24:0] n9401_o;
  wire [24:0] n9402_o;
  wire [24:0] n9403_o;
  wire [24:0] n9404_o;
  wire [24:0] n9405_o;
  wire n9407_o;
  wire [24:0] n9408_o;
  wire [24:0] n9409_o;
  wire [24:0] n9410_o;
  wire [24:0] n9411_o;
  wire [24:0] n9412_o;
  wire n9414_o;
  wire [24:0] n9415_o;
  wire [24:0] n9416_o;
  wire [24:0] n9417_o;
  wire [24:0] n9418_o;
  wire [24:0] n9419_o;
  wire n9421_o;
  wire [23:0] n9422_o;
  wire [23:0] n9423_o;
  wire [23:0] n9424_o;
  wire [23:0] n9425_o;
  wire [23:0] n9426_o;
  wire n9428_o;
  wire [15:0] n9429_o;
  wire [15:0] n9430_o;
  wire [15:0] n9431_o;
  wire [15:0] n9432_o;
  wire [15:0] n9433_o;
  wire n9435_o;
  wire [775:0] n9436_o;
  wire n9437_o;
  wire [775:0] n9438_o;
  wire [775:0] n9439_o;
  wire n9443_o;
  wire [31:0] n9444_o;
  wire [31:0] n9445_o;
  wire n9447_o;
  wire [31:0] n9448_o;
  wire [31:0] n9449_o;
  wire n9451_o;
  wire n9452_o;
  wire [63:0] n9454_o;
  wire n9456_o;
  wire n9457_o;
  wire [775:0] n9458_o;
  wire n9463_o;
  localparam [15:0] n9499_o = 16'bX;
  reg [15:0] n9498_source_is_safe_v;
  localparam [15:0] n9500_o = 16'bX;
  reg [15:0] n9498_dest_is_safe_v;
  wire n9502_o;
  wire n9504_o;
  wire n9505_o;
  wire n9506_o;
  wire n9507_o;
  wire n9508_o;
  wire n9509_o;
  wire n9510_o;
  wire n9511_o;
  wire n9512_o;
  wire n9513_o;
  wire n9514_o;
  wire n9515_o;
  wire n9516_o;
  wire n9517_o;
  wire n9518_o;
  wire n9519_o;
  wire n9520_o;
  wire n9521_o;
  wire n9522_o;
  wire n9523_o;
  wire n9524_o;
  wire n9525_o;
  wire n9526_o;
  wire n9527_o;
  wire n9528_o;
  wire n9529_o;
  wire n9530_o;
  wire n9531_o;
  wire n9532_o;
  wire n9533_o;
  wire n9534_o;
  wire n9535_o;
  wire n9536_o;
  wire n9537_o;
  wire n9538_o;
  wire n9539_o;
  wire n9540_o;
  wire n9541_o;
  wire n9542_o;
  wire n9543_o;
  wire n9544_o;
  wire n9545_o;
  wire n9546_o;
  wire n9547_o;
  wire n9548_o;
  wire n9549_o;
  wire n9550_o;
  wire n9551_o;
  wire n9552_o;
  wire n9553_o;
  wire n9554_o;
  wire n9555_o;
  wire n9556_o;
  wire n9557_o;
  wire n9558_o;
  wire n9559_o;
  wire n9560_o;
  wire n9561_o;
  wire n9562_o;
  wire n9563_o;
  wire n9564_o;
  wire n9565_o;
  wire n9566_o;
  wire n9567_o;
  wire n9568_o;
  wire n9569_o;
  wire n9570_o;
  wire n9571_o;
  wire n9572_o;
  wire n9573_o;
  wire n9574_o;
  wire n9575_o;
  wire n9576_o;
  wire n9577_o;
  wire n9578_o;
  wire n9579_o;
  wire n9580_o;
  wire n9581_o;
  wire n9582_o;
  wire n9583_o;
  wire n9584_o;
  wire n9585_o;
  wire n9586_o;
  wire n9587_o;
  wire n9588_o;
  wire n9589_o;
  wire n9590_o;
  wire n9591_o;
  wire n9592_o;
  wire n9593_o;
  wire n9594_o;
  wire n9595_o;
  wire [4:0] n9596_o;
  wire [15:0] n9597_o;
  wire n9598_o;
  wire n9599_o;
  wire n9600_o;
  wire [4:0] n9601_o;
  wire [15:0] n9602_o;
  wire n9603_o;
  wire n9604_o;
  wire n9605_o;
  wire n9606_o;
  wire [4:0] n9607_o;
  wire [15:0] n9608_o;
  wire n9609_o;
  wire n9610_o;
  wire n9611_o;
  wire [4:0] n9612_o;
  wire [15:0] n9613_o;
  wire n9614_o;
  wire n9615_o;
  wire n9616_o;
  wire n9617_o;
  wire [4:0] n9618_o;
  wire [15:0] n9619_o;
  wire n9620_o;
  wire n9621_o;
  wire n9622_o;
  wire [4:0] n9623_o;
  wire [15:0] n9624_o;
  wire n9625_o;
  wire n9626_o;
  wire n9627_o;
  wire n9628_o;
  wire [4:0] n9629_o;
  wire [15:0] n9630_o;
  wire n9631_o;
  wire n9632_o;
  wire n9633_o;
  wire [4:0] n9634_o;
  wire [15:0] n9635_o;
  wire n9636_o;
  wire n9637_o;
  wire n9638_o;
  wire n9639_o;
  wire [4:0] n9640_o;
  wire [15:0] n9641_o;
  wire n9642_o;
  wire n9643_o;
  wire n9644_o;
  wire [4:0] n9645_o;
  wire [15:0] n9646_o;
  wire n9647_o;
  wire n9648_o;
  wire n9649_o;
  wire n9650_o;
  wire [4:0] n9651_o;
  wire [15:0] n9652_o;
  wire n9653_o;
  wire n9654_o;
  wire n9655_o;
  wire [4:0] n9656_o;
  wire [15:0] n9657_o;
  wire n9658_o;
  wire n9659_o;
  wire n9660_o;
  wire n9661_o;
  wire [4:0] n9662_o;
  wire [15:0] n9663_o;
  wire n9664_o;
  wire n9665_o;
  wire n9666_o;
  wire [4:0] n9667_o;
  wire [15:0] n9668_o;
  wire n9669_o;
  wire n9670_o;
  wire n9671_o;
  wire n9672_o;
  wire [4:0] n9673_o;
  wire [15:0] n9674_o;
  wire n9675_o;
  wire n9676_o;
  wire n9677_o;
  wire [4:0] n9678_o;
  wire [15:0] n9679_o;
  wire n9680_o;
  wire n9681_o;
  wire n9682_o;
  wire n9683_o;
  wire [4:0] n9684_o;
  wire [15:0] n9685_o;
  wire n9686_o;
  wire n9687_o;
  wire n9688_o;
  wire [4:0] n9689_o;
  wire [15:0] n9690_o;
  wire n9691_o;
  wire n9692_o;
  wire [2:0] n9693_o;
  wire [2:0] n9694_o;
  wire [2:0] n9695_o;
  wire [2:0] n9702_o;
  wire [2:0] n9703_o;
  wire [2:0] n9704_o;
  wire [2:0] n9711_o;
  wire [2:0] n9712_o;
  wire [2:0] n9713_o;
  wire n9723_o;
  wire n9724_o;
  wire n9728_o;
  wire n9729_o;
  wire [4:0] n9733_o;
  wire [4:0] n9734_o;
  wire [2:0] n9748_o;
  wire n9749_o;
  wire [2:0] n9750_o;
  wire [2:0] n9751_o;
  reg [2:0] n9752_q;
  wire [2:0] n9753_o;
  wire n9754_o;
  wire [2:0] n9755_o;
  wire [2:0] n9756_o;
  reg [2:0] n9757_q;
  wire [2:0] n9758_o;
  wire n9759_o;
  wire [2:0] n9760_o;
  wire [2:0] n9761_o;
  reg [2:0] n9762_q;
  wire [15:0] n9766_o;
  wire [2:0] n9767_o;
  wire n9768_o;
  wire [2:0] n9769_o;
  wire [2:0] n9770_o;
  reg [2:0] n9771_q;
  wire [2:0] n9772_o;
  wire n9773_o;
  wire [2:0] n9774_o;
  wire [2:0] n9775_o;
  reg [2:0] n9776_q;
  wire [2:0] n9777_o;
  wire n9778_o;
  wire [2:0] n9779_o;
  wire [2:0] n9780_o;
  reg [2:0] n9781_q;
  wire [15:0] n9785_o;
  wire [1619:0] n9787_o;
  wire [2:0] n9788_o;
  wire n9790_o;
  wire [1619:0] n9791_o;
  wire [2:0] n9792_o;
  wire n9794_o;
  wire n9795_o;
  wire [1619:0] n9796_o;
  wire [3:0] n9797_o;
  wire n9799_o;
  wire n9800_o;
  wire [1619:0] n9801_o;
  wire n9802_o;
  wire [1619:0] n9803_o;
  wire n9804_o;
  wire n9805_o;
  wire n9806_o;
  wire n9807_o;
  wire [1619:0] n9808_o;
  wire [1:0] n9809_o;
  wire n9811_o;
  wire [1619:0] n9812_o;
  wire [1:0] n9813_o;
  wire n9815_o;
  wire n9816_o;
  wire n9817_o;
  wire n9818_o;
  wire n9819_o;
  wire [1619:0] n9820_o;
  wire [1:0] n9821_o;
  wire n9823_o;
  wire [1619:0] n9824_o;
  wire [1:0] n9825_o;
  wire n9827_o;
  wire n9828_o;
  wire n9829_o;
  wire n9830_o;
  wire n9831_o;
  wire n9832_o;
  wire [1619:0] n9833_o;
  wire [1:0] n9834_o;
  wire n9836_o;
  wire [1619:0] n9837_o;
  wire [1:0] n9838_o;
  wire n9840_o;
  wire n9841_o;
  wire n9842_o;
  wire n9843_o;
  wire n9844_o;
  wire n9845_o;
  wire n9846_o;
  wire n9851_o;
  wire n9852_o;
  wire [1619:0] n9853_o;
  wire n9854_o;
  wire n9856_o;
  wire n9857_o;
  wire n9858_o;
  wire n9859_o;
  wire [1619:0] n9860_o;
  wire n9861_o;
  wire n9863_o;
  wire [1619:0] n9864_o;
  wire n9865_o;
  wire n9867_o;
  wire [1619:0] n9868_o;
  wire [1:0] n9869_o;
  wire [1:0] n9870_o;
  wire [1:0] n9871_o;
  wire n9872_o;
  wire n9873_o;
  wire [1619:0] n9874_o;
  wire [1:0] n9875_o;
  wire [1:0] n9876_o;
  wire n9877_o;
  wire n9878_o;
  wire n9883_o;
  wire [1619:0] n9885_o;
  wire [2:0] n9886_o;
  wire n9888_o;
  wire [1619:0] n9889_o;
  wire [3:0] n9890_o;
  wire [3:0] n9891_o;
  wire [3:0] n9892_o;
  wire n9894_o;
  wire n9895_o;
  wire [1619:0] n9897_o;
  wire [2:0] n9898_o;
  wire n9900_o;
  wire [1619:0] n9901_o;
  wire n9902_o;
  wire n9903_o;
  wire n9904_o;
  wire [1619:0] n9905_o;
  wire [3:0] n9906_o;
  wire [3:0] n9907_o;
  wire n9909_o;
  wire n9910_o;
  wire [1619:0] n9912_o;
  wire [2:0] n9913_o;
  wire n9915_o;
  wire [1619:0] n9916_o;
  wire n9917_o;
  wire n9918_o;
  wire [1619:0] n9919_o;
  wire [3:0] n9920_o;
  wire [3:0] n9921_o;
  wire n9923_o;
  wire n9924_o;
  wire [1619:0] n9926_o;
  wire [2:0] n9927_o;
  wire n9929_o;
  wire [1619:0] n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9933_o;
  wire n9936_o;
  wire [1619:0] n9937_o;
  wire [2:0] n9938_o;
  wire n9940_o;
  wire [1619:0] n9941_o;
  wire n9942_o;
  wire n9943_o;
  wire n9946_o;
  wire [1619:0] n9947_o;
  wire [2:0] n9948_o;
  wire n9950_o;
  wire [1619:0] n9951_o;
  wire [1:0] n9952_o;
  wire n9954_o;
  wire [1619:0] n9955_o;
  wire n9956_o;
  wire n9957_o;
  wire n9958_o;
  wire [1619:0] n9959_o;
  wire [1:0] n9960_o;
  wire n9962_o;
  wire [1619:0] n9963_o;
  wire n9964_o;
  wire n9965_o;
  wire n9966_o;
  wire n9967_o;
  wire n9968_o;
  wire [1619:0] n9970_o;
  wire [1:0] n9971_o;
  wire [1619:0] n9974_o;
  wire [1:0] n9975_o;
  wire n9980_o;
  wire n9981_o;
  wire n9983_o;
  wire n9984_o;
  wire n9985_o;
  wire n9986_o;
  wire n9987_o;
  wire n9988_o;
  wire n9989_o;
  wire n9991_o;
  wire n9992_o;
  wire [1619:0] n9994_o;
  wire [2:0] n9995_o;
  wire n9997_o;
  wire [1619:0] n9998_o;
  wire [3:0] n9999_o;
  wire [3:0] n10000_o;
  wire [3:0] n10001_o;
  wire n10003_o;
  wire n10004_o;
  wire [1619:0] n10006_o;
  wire [2:0] n10007_o;
  wire n10009_o;
  wire [1619:0] n10010_o;
  wire n10011_o;
  wire n10012_o;
  wire n10013_o;
  wire [1619:0] n10014_o;
  wire [3:0] n10015_o;
  wire [3:0] n10016_o;
  wire n10018_o;
  wire n10019_o;
  wire [1619:0] n10021_o;
  wire [2:0] n10022_o;
  wire n10024_o;
  wire [1619:0] n10025_o;
  wire n10026_o;
  wire n10027_o;
  wire [1619:0] n10028_o;
  wire [3:0] n10029_o;
  wire [3:0] n10030_o;
  wire n10032_o;
  wire n10033_o;
  wire [1619:0] n10035_o;
  wire [2:0] n10036_o;
  wire n10038_o;
  wire [1619:0] n10039_o;
  wire n10040_o;
  wire n10041_o;
  wire n10042_o;
  wire n10045_o;
  wire [1619:0] n10046_o;
  wire [2:0] n10047_o;
  wire n10049_o;
  wire [1619:0] n10050_o;
  wire n10051_o;
  wire n10052_o;
  wire n10055_o;
  wire [1619:0] n10056_o;
  wire [2:0] n10057_o;
  wire n10059_o;
  wire [1619:0] n10060_o;
  wire [1:0] n10061_o;
  wire n10063_o;
  wire [1619:0] n10064_o;
  wire n10065_o;
  wire n10066_o;
  wire n10067_o;
  wire [1619:0] n10068_o;
  wire [1:0] n10069_o;
  wire n10071_o;
  wire [1619:0] n10072_o;
  wire n10073_o;
  wire n10074_o;
  wire n10075_o;
  wire n10076_o;
  wire n10077_o;
  wire [1619:0] n10079_o;
  wire [1:0] n10080_o;
  wire [1619:0] n10083_o;
  wire [1:0] n10084_o;
  wire n10089_o;
  wire n10090_o;
  wire n10092_o;
  wire n10093_o;
  wire n10094_o;
  wire n10095_o;
  wire n10096_o;
  wire n10097_o;
  wire n10098_o;
  wire n10100_o;
  wire [2:0] n10104_o;
  wire n10106_o;
  wire n10107_o;
  wire n10108_o;
  wire n10109_o;
  wire n10112_o;
  wire n10116_o;
  wire [63:0] n10118_o;
  wire [2:0] n10119_o;
  wire n10121_o;
  wire n10122_o;
  wire n10123_o;
  wire n10124_o;
  wire n10127_o;
  wire [2:0] n10144_o;
  wire n10146_o;
  wire n10147_o;
  wire n10148_o;
  wire n10149_o;
  wire n10150_o;
  wire n10151_o;
  wire n10152_o;
  wire [10:0] n10153_o;
  wire [4:0] n10154_o;
  wire n10155_o;
  wire [1:0] n10156_o;
  wire [3:0] n10157_o;
  wire [1:0] n10158_o;
  wire [12:0] n10159_o;
  wire [12:0] n10160_o;
  wire [2:0] n10161_o;
  wire n10163_o;
  wire n10164_o;
  wire n10165_o;
  wire n10166_o;
  wire n10167_o;
  wire n10168_o;
  wire [10:0] n10169_o;
  wire [4:0] n10170_o;
  wire n10171_o;
  wire [1:0] n10172_o;
  wire [3:0] n10173_o;
  wire [1:0] n10174_o;
  wire [12:0] n10175_o;
  wire [12:0] n10176_o;
  wire [10:0] n10178_o;
  wire [4:0] n10180_o;
  wire [3:0] n10182_o;
  wire [1:0] n10184_o;
  wire [27:0] n10185_o;
  wire [27:0] n10187_o;
  wire n10189_o;
  wire n10192_o;
  wire n10195_o;
  wire [10:0] n10198_o;
  wire [4:0] n10199_o;
  wire [3:0] n10200_o;
  wire [1:0] n10201_o;
  wire [27:0] n10202_o;
  wire [27:0] n10203_o;
  wire n10204_o;
  wire n10206_o;
  wire n10208_o;
  wire [2:0] n10214_o;
  wire n10216_o;
  wire n10217_o;
  wire n10219_o;
  wire n10221_o;
  wire n10225_o;
  wire n10227_o;
  wire n10228_o;
  wire [2:0] n10229_o;
  wire n10231_o;
  wire [2:0] n10232_o;
  wire n10234_o;
  wire n10236_o;
  wire n10238_o;
  wire n10246_o;
  wire n10248_o;
  wire n10250_o;
  wire n10258_o;
  wire n10292_o;
  wire n10294_o;
  wire n10295_o;
  wire [1:0] n10297_o;
  wire n10298_o;
  wire [1:0] n10299_o;
  wire [1:0] n10301_o;
  wire n10302_o;
  wire [1:0] n10303_o;
  wire [1:0] n10304_o;
  wire [1:0] n10305_o;
  wire [1:0] n10306_o;
  wire [1:0] n10307_o;
  wire [1:0] n10308_o;
  wire [1:0] n10309_o;
  wire [1:0] n10310_o;
  wire n10311_o;
  wire n10312_o;
  wire n10313_o;
  wire n10314_o;
  wire [1:0] n10315_o;
  wire [1:0] n10316_o;
  wire [1:0] n10317_o;
  wire [1:0] n10318_o;
  wire [1:0] n10320_o;
  wire [3:0] n10321_o;
  wire [3:0] n10322_o;
  wire [1:0] n10323_o;
  wire [1:0] n10324_o;
  wire [3:0] n10325_o;
  wire [3:0] n10326_o;
  wire n10356_o;
  wire n10359_o;
  wire n10362_o;
  wire [23:0] n10363_o;
  wire [23:0] n10364_o;
  wire n10365_o;
  wire n10368_o;
  wire [23:0] n10369_o;
  wire [23:0] n10370_o;
  wire n10371_o;
  wire n10374_o;
  wire [23:0] n10375_o;
  wire [23:0] n10376_o;
  wire n10377_o;
  wire n10380_o;
  wire [23:0] n10381_o;
  wire [23:0] n10382_o;
  wire n10383_o;
  wire n10386_o;
  wire n10387_o;
  wire n10390_o;
  wire n10392_o;
  wire [23:0] n10393_o;
  wire [775:0] n10394_o;
  wire n10395_o;
  wire [1:0] n10396_o;
  wire n10398_o;
  wire n10399_o;
  wire [23:0] n10401_o;
  wire [23:0] n10402_o;
  wire [1:0] n10403_o;
  wire n10405_o;
  wire n10406_o;
  wire n10407_o;
  wire [23:0] n10408_o;
  wire [23:0] n10409_o;
  wire [23:0] n10411_o;
  wire [23:0] n10412_o;
  wire [23:0] n10414_o;
  wire [23:0] n10415_o;
  wire [23:0] n10416_o;
  wire [23:0] n10417_o;
  wire n10418_o;
  wire n10419_o;
  wire [1:0] n10420_o;
  wire n10422_o;
  wire n10423_o;
  wire n10424_o;
  wire [23:0] n10425_o;
  wire [23:0] n10426_o;
  wire [23:0] n10428_o;
  wire [23:0] n10429_o;
  wire [23:0] n10431_o;
  wire [23:0] n10432_o;
  wire [23:0] n10433_o;
  wire [23:0] n10434_o;
  wire n10435_o;
  wire n10436_o;
  wire [23:0] n10437_o;
  wire [47:0] n10438_o;
  wire [47:0] n10439_o;
  wire [23:0] n10440_o;
  wire [1:0] n10441_o;
  wire [1:0] n10442_o;
  wire [1:0] n10443_o;
  wire n10445_o;
  wire [47:0] n10446_o;
  wire [47:0] n10448_o;
  wire [23:0] n10449_o;
  wire [1:0] n10450_o;
  wire [1:0] n10451_o;
  wire [1:0] n10452_o;
  wire [1:0] n10453_o;
  wire [1:0] n10454_o;
  wire n10455_o;
  wire n10456_o;
  wire [1:0] n10459_o;
  wire [1:0] n10460_o;
  wire [1:0] n10461_o;
  wire [1:0] n10462_o;
  wire n10463_o;
  wire n10466_o;
  wire [1:0] n10467_o;
  wire n10469_o;
  wire n10470_o;
  wire n10471_o;
  wire n10472_o;
  wire n10473_o;
  wire n10476_o;
  wire [1:0] n10477_o;
  wire n10479_o;
  wire n10480_o;
  wire n10481_o;
  wire n10482_o;
  wire n10483_o;
  wire n10485_o;
  wire n10486_o;
  wire n10489_o;
  wire n10490_o;
  wire n10491_o;
  wire n10493_o;
  wire [1:0] n10494_o;
  wire n10496_o;
  wire n10497_o;
  wire n10498_o;
  wire n10499_o;
  wire n10502_o;
  wire [1:0] n10503_o;
  wire n10505_o;
  wire n10506_o;
  wire n10507_o;
  wire n10508_o;
  wire n10510_o;
  wire n10511_o;
  wire n10514_o;
  wire n10515_o;
  wire n10516_o;
  wire n10518_o;
  wire [1:0] n10519_o;
  wire n10521_o;
  wire n10522_o;
  wire n10523_o;
  wire n10524_o;
  wire n10525_o;
  wire n10528_o;
  wire [1:0] n10529_o;
  wire n10531_o;
  wire n10532_o;
  wire n10533_o;
  wire n10534_o;
  wire n10535_o;
  wire n10537_o;
  wire n10538_o;
  wire n10541_o;
  wire n10542_o;
  wire n10543_o;
  wire n10545_o;
  wire [1:0] n10546_o;
  wire n10548_o;
  wire n10549_o;
  wire n10550_o;
  wire n10551_o;
  wire n10554_o;
  wire [1:0] n10555_o;
  wire n10557_o;
  wire n10558_o;
  wire n10559_o;
  wire n10560_o;
  wire n10562_o;
  wire n10563_o;
  wire n10566_o;
  wire n10567_o;
  wire n10568_o;
  wire n10570_o;
  wire [1:0] n10571_o;
  wire n10573_o;
  wire n10574_o;
  wire n10576_o;
  wire [1:0] n10577_o;
  wire n10579_o;
  wire n10580_o;
  wire n10581_o;
  wire n10582_o;
  wire n10583_o;
  wire n10586_o;
  wire n10588_o;
  wire n10590_o;
  wire [1:0] n10591_o;
  wire n10593_o;
  wire n10594_o;
  wire n10595_o;
  wire n10596_o;
  wire n10597_o;
  wire n10598_o;
  wire n10599_o;
  wire [1:0] n10600_o;
  wire n10602_o;
  wire n10603_o;
  wire n10604_o;
  wire n10605_o;
  wire n10606_o;
  wire n10607_o;
  wire n10608_o;
  wire n10609_o;
  wire n10610_o;
  wire n10611_o;
  wire n10612_o;
  wire n10613_o;
  wire n10614_o;
  wire n10615_o;
  wire n10618_o;
  wire [1:0] n10619_o;
  wire n10621_o;
  wire n10622_o;
  wire n10623_o;
  wire n10624_o;
  wire n10625_o;
  wire n10626_o;
  wire [1:0] n10627_o;
  wire n10629_o;
  wire n10630_o;
  wire n10631_o;
  wire n10632_o;
  wire n10633_o;
  wire n10634_o;
  wire n10635_o;
  wire n10636_o;
  wire n10637_o;
  wire n10638_o;
  wire n10639_o;
  wire n10640_o;
  wire n10641_o;
  wire n10644_o;
  wire [1:0] n10645_o;
  wire n10647_o;
  wire n10648_o;
  wire n10649_o;
  wire n10650_o;
  wire n10651_o;
  wire n10652_o;
  wire n10653_o;
  wire [1:0] n10654_o;
  wire n10656_o;
  wire n10657_o;
  wire n10658_o;
  wire n10659_o;
  wire n10660_o;
  wire n10661_o;
  wire n10662_o;
  wire n10663_o;
  wire n10664_o;
  wire n10665_o;
  wire n10666_o;
  wire n10667_o;
  wire n10668_o;
  wire n10669_o;
  wire n10672_o;
  wire [1:0] n10673_o;
  wire n10675_o;
  wire n10676_o;
  wire n10677_o;
  wire n10678_o;
  wire n10679_o;
  wire n10680_o;
  wire [1:0] n10681_o;
  wire n10683_o;
  wire n10684_o;
  wire n10685_o;
  wire n10686_o;
  wire n10687_o;
  wire n10688_o;
  wire n10689_o;
  wire n10690_o;
  wire n10691_o;
  wire n10692_o;
  wire n10693_o;
  wire n10694_o;
  wire n10695_o;
  wire n10698_o;
  wire [1:0] n10699_o;
  wire n10701_o;
  wire n10702_o;
  wire n10703_o;
  wire n10704_o;
  wire [1:0] n10705_o;
  wire n10707_o;
  wire n10708_o;
  wire n10709_o;
  wire n10710_o;
  wire n10711_o;
  wire n10712_o;
  wire n10713_o;
  wire n10714_o;
  wire n10715_o;
  wire n10716_o;
  wire n10717_o;
  wire n10720_o;
  wire n10722_o;
  wire [1:0] n10723_o;
  wire n10725_o;
  wire n10726_o;
  wire n10727_o;
  wire n10728_o;
  wire n10729_o;
  wire n10731_o;
  wire n10733_o;
  wire [1:0] n10734_o;
  wire n10736_o;
  wire n10737_o;
  wire n10738_o;
  wire n10739_o;
  wire n10741_o;
  wire n10743_o;
  wire [1:0] n10744_o;
  wire n10746_o;
  wire n10747_o;
  wire n10748_o;
  wire n10749_o;
  wire n10750_o;
  wire n10752_o;
  wire n10754_o;
  wire [1:0] n10755_o;
  wire n10757_o;
  wire n10758_o;
  wire n10759_o;
  wire n10760_o;
  wire n10762_o;
  wire n10764_o;
  wire [1:0] n10765_o;
  wire n10767_o;
  wire n10768_o;
  wire n10770_o;
  wire [1:0] n10771_o;
  wire n10772_o;
  wire [1:0] n10773_o;
  wire n10774_o;
  wire n10775_o;
  wire [1:0] n10776_o;
  wire n10777_o;
  wire [1:0] n10778_o;
  wire n10779_o;
  wire n10780_o;
  wire n10781_o;
  wire [1:0] n10782_o;
  wire n10783_o;
  wire [1:0] n10784_o;
  wire n10785_o;
  wire n10786_o;
  wire [1:0] n10787_o;
  wire n10788_o;
  wire [1:0] n10789_o;
  wire n10790_o;
  wire n10791_o;
  wire n10792_o;
  wire [1:0] n10793_o;
  wire n10794_o;
  wire [1:0] n10795_o;
  wire n10796_o;
  wire [1:0] n10797_o;
  wire [1:0] n10798_o;
  wire [1:0] n10799_o;
  wire [1:0] n10803_o;
  wire [1:0] n10811_o;
  wire [1:0] n10816_o;
  wire n10858_o;
  wire n10859_o;
  wire n10865_o;
  wire n10866_o;
  wire n10908_o;
  wire [31:0] n10911_o;
  wire [1:0] n10912_o;
  wire n10914_o;
  wire n10915_o;
  wire [3239:0] n10924_o;
  wire [1:0] n10925_o;
  wire [1:0] n10926_o;
  wire [47:0] n10927_o;
  reg [47:0] n10928_q;
  wire [47:0] n10929_o;
  reg [47:0] n10930_q;
  wire [23:0] n10931_o;
  reg [23:0] n10932_q;
  reg [1:0] n10933_q;
  reg [1:0] n10934_q;
  reg n10935_q;
  reg [1:0] n10936_q;
  reg [1:0] n10937_q;
  reg n10938_q;
  wire n10939_o;
  reg n10940_q;
  reg n10941_q;
  reg n10942_q;
  reg [63:0] n10943_q;
  reg [63:0] n10944_q;
  reg n10945_q;
  wire [63:0] n10946_o;
  reg [63:0] n10947_q;
  wire [31:0] n10948_o;
  reg [31:0] n10949_q;
  wire n10950_o;
  reg n10951_q;
  wire [31:0] n10952_o;
  reg [31:0] n10953_q;
  reg [1:0] n10954_q;
  reg [1:0] n10955_q;
  wire n10956_o;
  wire [1619:0] n10957_o;
  reg [1619:0] n10958_q;
  wire n10959_o;
  wire [1619:0] n10960_o;
  reg [1619:0] n10961_q;
  wire [63:0] n10962_o;
  reg [63:0] n10963_q;
  wire [31:0] n10964_o;
  reg [31:0] n10965_q;
  reg [31:0] n10966_q;
  reg n10968_q;
  wire [3:0] n10969_o;
  reg [3:0] n10970_q;
  reg [3:0] n10971_q;
  reg [1:0] n10972_q;
  reg [3:0] n10973_q;
  reg [2:0] n10974_q;
  reg [2:0] n10975_q;
  reg [2:0] n10976_q;
  wire [15:0] n10977_o;
  reg n10978_q;
  reg [1:0] n10979_q;
  wire [3:0] n10980_o;
  reg n10981_q;
  reg [1:0] n10982_q;
  wire [3:0] n10983_o;
  wire n10984_o;
  reg n10985_q;
  reg [1:0] n10986_q;
  reg [1:0] n10987_q;
  reg n10988_q;
  wire [775:0] n10989_o;
  reg [775:0] n10990_q;
  wire [775:0] n10991_o;
  reg [775:0] n10992_q;
  reg [775:0] n10993_q;
  wire [1:0] n10994_o;
  wire [10:0] n10995_o;
  reg [10:0] n10996_q;
  wire [4:0] n10997_o;
  reg [4:0] n10998_q;
  wire [3:0] n10999_o;
  reg [3:0] n11000_q;
  wire [1:0] n11001_o;
  reg [1:0] n11002_q;
  wire [27:0] n11003_o;
  reg [27:0] n11004_q;
  wire n11005_o;
  reg n11006_q;
  reg n11007_q;
  wire n11008_o;
  reg n11009_q;
  reg [11:0] n11011_q;
  reg [11:0] n11012_q;
  reg n11013_q;
  reg n11014_q;
  reg [31:0] n11015_q;
  reg n11016_q;
  wire n11017_o;
  wire n11018_o;
  wire n11019_o;
  wire n11020_o;
  wire n11021_o;
  wire n11022_o;
  wire n11023_o;
  wire n11024_o;
  wire n11025_o;
  wire n11026_o;
  wire n11027_o;
  wire n11028_o;
  wire n11029_o;
  wire n11030_o;
  wire n11031_o;
  wire n11032_o;
  wire [3:0] n11033_o;
  wire [1:0] n11034_o;
  reg n11035_o;
  wire [1:0] n11036_o;
  reg n11037_o;
  wire [1:0] n11038_o;
  reg n11039_o;
  wire [1:0] n11040_o;
  reg n11041_o;
  wire [1:0] n11042_o;
  reg n11043_o;
  wire n11044_o;
  wire n11045_o;
  wire n11046_o;
  wire n11047_o;
  wire n11048_o;
  wire n11049_o;
  wire n11050_o;
  wire n11051_o;
  wire n11052_o;
  wire n11053_o;
  wire n11054_o;
  wire n11055_o;
  wire n11056_o;
  wire n11057_o;
  wire n11058_o;
  wire n11059_o;
  wire [3:0] n11060_o;
  wire [1:0] n11061_o;
  reg n11062_o;
  wire [1:0] n11063_o;
  reg n11064_o;
  wire [1:0] n11065_o;
  reg n11066_o;
  wire [1:0] n11067_o;
  reg n11068_o;
  wire [1:0] n11069_o;
  reg n11070_o;
  assign bus_readdata_out = bus_readdata_r;
  assign bus_readdatavalid_out = rden_r;
  assign bus_writewait_out = waitrequest;
  assign bus_readwait_out = n7857_o;
  assign instruction_valid_out = instruction_valid_rr;
  assign instruction_out_opcode = n7776_o;
  assign instruction_out_condition = n7777_o;
  assign instruction_out_vm = n7778_o;
  assign instruction_out_source = n7779_o;
  assign instruction_out_source_bus_id = n7780_o;
  assign instruction_out_source_data_type = n7781_o;
  assign instruction_out_dest = n7782_o;
  assign instruction_out_dest_bus_id = n7783_o;
  assign instruction_out_dest_data_type = n7784_o;
  assign instruction_out_mcast = n7785_o;
  assign instruction_out_count = n7786_o;
  assign instruction_out_data = n7787_o;
  assign instruction_out_repeat = n7788_o;
  assign instruction_out_source_addr_mode = n7789_o;
  assign instruction_out_dest_addr_mode = n7790_o;
  assign instruction_out_stream_process = n7791_o;
  assign instruction_out_stream_process_id = n7792_o;
  assign pre_instruction_out_opcode = n7794_o;
  assign pre_instruction_out_condition = n7795_o;
  assign pre_instruction_out_vm = n7796_o;
  assign pre_instruction_out_source = n7797_o;
  assign pre_instruction_out_source_bus_id = n7798_o;
  assign pre_instruction_out_source_data_type = n7799_o;
  assign pre_instruction_out_dest = n7800_o;
  assign pre_instruction_out_dest_bus_id = n7801_o;
  assign pre_instruction_out_dest_data_type = n7802_o;
  assign pre_instruction_out_mcast = n7803_o;
  assign pre_instruction_out_count = n7804_o;
  assign pre_instruction_out_data = n7805_o;
  assign pre_instruction_out_repeat = n7806_o;
  assign pre_instruction_out_source_addr_mode = n7807_o;
  assign pre_instruction_out_dest_addr_mode = n7808_o;
  assign pre_instruction_out_stream_process = n7809_o;
  assign pre_instruction_out_stream_process_id = n7810_o;
  assign task_start_addr_out = task_start_addr_r;
  assign task_pending_out = task_r;
  assign task_out = task2;
  assign task_vm_out = task_vm_r;
  assign task_pcore_out = task_pcore_r;
  assign task_lockstep_out = task_lockstep_r;
  assign task_tid_mask_out = task_tid_mask_r;
  assign task_iregister_auto_out = task_iregister_auto_r;
  assign task_data_model_out = task_data_model_r;
  assign indication_avail_out = n7826_o;
  /* ../../HW/platform/simulation/DPRAM.vhd:42:9  */
  assign n7776_o = instruction_rr[2:0];
  /* ../../HW/src/top/cell.vhd:166:10  */
  assign n7777_o = instruction_rr[6:3];
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  assign n7778_o = instruction_rr[7];
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
  assign n7779_o = instruction_rr[783:8];
  /* ../../HW/platform/simulation/DPRAM.vhd:58:1  */
  assign n7780_o = instruction_rr[785:784];
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  assign n7781_o = instruction_rr[787:786];
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  assign n7782_o = instruction_rr[1563:788];
  /* ../../HW/src/top/cell.vhd:165:10  */
  assign n7783_o = instruction_rr[1565:1564];
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign n7784_o = instruction_rr[1567:1566];
  /* ../../HW/src/top/cell.vhd:164:10  */
  assign n7785_o = instruction_rr[1573:1568];
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign n7786_o = instruction_rr[1597:1574];
  /* ../../HW/src/top/cell.vhd:163:10  */
  assign n7787_o = instruction_rr[1613:1598];
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign n7788_o = instruction_rr[1614];
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7789_o = instruction_rr[1615];
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign n7790_o = instruction_rr[1616];
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7791_o = instruction_rr[1617];
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7792_o = instruction_rr[1619:1618];
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign n7794_o = instruction_r[2:0];
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7795_o = instruction_r[6:3];
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7796_o = instruction_r[7];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7797_o = instruction_r[783:8];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7798_o = instruction_r[785:784];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7799_o = instruction_r[787:786];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7800_o = instruction_r[1563:788];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7801_o = instruction_r[1565:1564];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7802_o = instruction_r[1567:1566];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7803_o = instruction_r[1573:1568];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7804_o = instruction_r[1597:1574];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7805_o = instruction_r[1613:1598];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7806_o = instruction_r[1614];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7807_o = instruction_r[1615];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7808_o = instruction_r[1616];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7809_o = instruction_r[1617];
  /* ../../HW/src/top/cell.vhd:322:1  */
  assign n7810_o = instruction_r[1619:1618];
  /* ../../HW/src/dp/dp_fetch.vhd:140:8  */
  assign fifo_avail = fifo_i_n7936; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:141:8  */
  assign match = 1'b1; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:142:8  */
  assign irec = n8819_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:143:8  */
  assign irec_generic = n8835_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:144:8  */
  assign orec = n9874_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:145:8  */
  assign orecs = n10924_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:146:8  */
  assign orec_generic = n8779_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:147:8  */
  assign data = n8398_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:148:8  */
  assign q1 = fifo_i_n7929; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:149:8  */
  assign q2 = fifo_i_n7930; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:150:8  */
  assign rdreq = n7927_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:151:8  */
  assign rdreqs = n9876_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:152:8  */
  assign wreq = n8842_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:153:8  */
  assign wreq_all = n8840_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:154:8  */
  assign full = fifo_i_n7935; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:155:8  */
  assign ready = n8900_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:156:8  */
  assign ready_which = n8902_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:157:8  */
  assign ready2 = n10925_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:158:8  */
  assign valid = n9877_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:159:8  */
  assign valids = n10926_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:160:8  */
  assign wregno = n8152_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:161:8  */
  assign rregno = n8155_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:162:8  */
  assign pcore_sink_counter_r = n10928_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:163:8  */
  assign sram_sink_counter_r = n10930_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:164:8  */
  assign ddr_sink_counter_r = n10932_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:165:8  */
  assign sink_pcore_busy_r = n10933_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:166:8  */
  assign sink_sram_busy_r = n10934_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:167:8  */
  assign sink_ddr_busy_r = n10935_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:168:8  */
  assign pcore_source_busy_r = n10936_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:169:8  */
  assign sram_source_busy_r = n10937_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:170:8  */
  assign ddr_source_busy_r = n10938_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:171:8  */
  assign log_enable_r = n10940_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:172:8  */
  assign print_indication_r = n10941_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:173:8  */
  assign print_indication_rr = n10942_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:174:8  */
  assign print_param_r = n10943_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:175:8  */
  assign print_param_rr = n10944_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:176:8  */
  assign wreq2 = n10221_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:177:8  */
  assign wreq2_indication = n10112_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:178:8  */
  assign pcore_read_pending = n8149_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:179:8  */
  assign sram_read_pending = n8150_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:180:8  */
  assign ddr_read_pending = n8151_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:186:8  */
  assign indication_full_r = n10945_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:188:8  */
  assign indication_rdreq = n8909_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:189:8  */
  assign in_indication = n8131_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:190:8  */
  assign indication = indication_i_n8132; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:191:8  */
  assign indication_rdusedw = indication_i_n8133; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:192:8  */
  assign indication_wrusedw = indication_i_n8134; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:193:8  */
  assign indication_parm_r = n10947_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:194:8  */
  assign indication_r = n10949_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:195:8  */
  assign indication_sync_r = n10951_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:199:8  */
  assign bus_readdata_r = n10953_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:201:8  */
  assign instruction_valid_r = n10954_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:202:8  */
  assign instruction_valid_rr = n10955_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:203:8  */
  assign instruction_r = n10958_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:204:8  */
  assign instruction_rr = n10961_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:205:8  */
  assign instruction = orec; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:207:8  */
  assign log_status_last_r = n10963_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:208:8  */
  assign log_write = n7901_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:209:8  */
  assign log_read = log_fifo_i_n7908; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:210:8  */
  assign log_readtime_r = n10965_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:211:8  */
  assign log_rdreq = n8918_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:212:8  */
  assign log_empty = log_fifo_i_n7911; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:213:8  */
  assign log_full = log_fifo_i_n7912; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:214:8  */
  assign log_time_r = n10966_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:216:8  */
  assign log_wrreq = n7903_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:217:8  */
  assign log_wrreq2 = n7907_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:219:8  */
  assign load = n7865_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:220:8  */
  assign load_r = n10968_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:221:8  */
  assign load_busid_r = n10970_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:223:8  */
  assign dp_var_waddress = load_busid_r; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:224:8  */
  assign dp_var_raddress = n8126_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:225:8  */
  assign dp_var_write = n8037_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:226:8  */
  assign dp_var_read = gen1_ram_i_n7949; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:227:8  */
  assign dp_var_we = load_r; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:228:8  */
  assign dp_var_template = n8123_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:230:8  */
  assign task2 = n7835_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:231:8  */
  assign waitrequest = n7855_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:235:8  */
  assign source_bus_id_r = n10971_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:236:8  */
  assign source_vm_r = n10972_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:237:8  */
  assign dest_bus_id_r = n10973_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:239:8  */
  assign outoforderok = n9846_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:243:8  */
  assign new_cmd_is_safe_r = n10977_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:244:8  */
  assign condition_vm0_busy_r = n10980_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:245:8  */
  assign condition_vm1_busy_r = n10983_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:247:8  */
  assign curr_vm_r = n10985_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:249:8  */
  assign pcore_sink_busy_r = n10986_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:250:8  */
  assign sram_sink_busy_r = n10987_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:251:8  */
  assign ddr_sink_busy_r = n10988_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:899:8  */
  assign wregno2 = n8153_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:901:8  */
  assign wregno2_r = n8154_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:903:8  */
  always @*
    src_template_r = n10990_q; // (isignal)
  initial
    src_template_r = 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:904:8  */
  always @*
    dest_template_r = n10992_q; // (isignal)
  initial
    dest_template_r = 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:905:8  */
  always @*
    template_r = n10993_q; // (isignal)
  initial
    template_r = 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:906:8  */
  assign pause = n9878_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:907:8  */
  assign pauses = n10994_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:908:8  */
  assign task_start_addr = n10198_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:909:8  */
  assign task_pcore = n10199_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:910:8  */
  assign task_tid_mask = n10200_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:911:8  */
  assign task_data_model = n10201_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:912:8  */
  assign task_iregister_auto = n10203_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:913:8  */
  assign task_lockstep = n10204_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:914:8  */
  assign \task  = n10206_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:915:8  */
  assign task_vm = n10208_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:916:8  */
  assign task_start_addr_r = n10996_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:917:8  */
  always @*
    task_pcore_r = n10998_q; // (isignal)
  initial
    task_pcore_r = 5'b11111;
  /* ../../HW/src/dp/dp_fetch.vhd:918:8  */
  always @*
    task_tid_mask_r = n11000_q; // (isignal)
  initial
    task_tid_mask_r = 4'b1111;
  /* ../../HW/src/dp/dp_fetch.vhd:919:8  */
  assign task_data_model_r = n11002_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:920:8  */
  assign task_iregister_auto_r = n11004_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:921:8  */
  assign task_lockstep_r = n11006_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:922:8  */
  assign task_r = n11007_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:923:8  */
  assign task_vm_r = n11009_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:925:8  */
  assign bus_waddr_r = n11011_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:926:8  */
  assign bus_raddr_r = n11012_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:927:8  */
  assign bus_write_r = n11013_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:928:8  */
  assign bus_read_r = n11014_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:929:8  */
  assign bus_writedata_r = n11015_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:930:8  */
  assign rden_r = n11016_q; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:931:8  */
  assign avail = n7846_o; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:932:8  */
  assign indication_empty = indication_i_n8135; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:935:25  */
  assign n7826_o = ~indication_empty;
  /* ../../HW/src/dp/dp_fetch.vhd:938:18  */
  assign n7827_o = task_r & task_ready_in;
  /* ../../HW/src/dp/dp_fetch.vhd:938:64  */
  assign n7828_o = pcore_source_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:938:41  */
  assign n7829_o = ~n7828_o;
  /* ../../HW/src/dp/dp_fetch.vhd:938:36  */
  assign n7830_o = n7827_o & n7829_o;
  /* ../../HW/src/dp/dp_fetch.vhd:938:95  */
  assign n7831_o = sink_pcore_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:938:74  */
  assign n7832_o = ~n7831_o;
  /* ../../HW/src/dp/dp_fetch.vhd:938:69  */
  assign n7833_o = n7830_o & n7832_o;
  /* ../../HW/src/dp/dp_fetch.vhd:938:115  */
  assign n7834_o = ~task_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:938:101  */
  assign n7835_o = n7834_o ? n7833_o : n7842_o;
  /* ../../HW/src/dp/dp_fetch.vhd:940:18  */
  assign n7836_o = task_r & task_ready_in;
  /* ../../HW/src/dp/dp_fetch.vhd:940:64  */
  assign n7837_o = pcore_source_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:940:41  */
  assign n7838_o = ~n7837_o;
  /* ../../HW/src/dp/dp_fetch.vhd:940:36  */
  assign n7839_o = n7836_o & n7838_o;
  /* ../../HW/src/dp/dp_fetch.vhd:940:95  */
  assign n7840_o = sink_pcore_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:940:74  */
  assign n7841_o = ~n7840_o;
  /* ../../HW/src/dp/dp_fetch.vhd:940:69  */
  assign n7842_o = n7839_o & n7841_o;
  /* ../../HW/src/dp/dp_fetch.vhd:949:24  */
  assign n7843_o = ~instruction_valid_r;
  /* ../../HW/src/dp/dp_fetch.vhd:949:19  */
  assign n7844_o = ready_in & n7843_o;
  /* ../../HW/src/dp/dp_fetch.vhd:949:54  */
  assign n7845_o = ~instruction_valid_rr;
  /* ../../HW/src/dp/dp_fetch.vhd:949:49  */
  assign n7846_o = n7844_o & n7845_o;
  /* ../../HW/src/dp/dp_fetch.vhd:953:36  */
  assign n7848_o = full | load;
  /* ../../HW/src/dp/dp_fetch.vhd:953:48  */
  assign n7849_o = n7848_o | wreq;
  /* ../../HW/src/dp/dp_fetch.vhd:953:86  */
  assign n7850_o = bus_waddr_in[4:0];
  /* ../../HW/src/dp/dp_fetch.vhd:953:117  */
  assign n7852_o = n7850_o == 5'b00101;
  /* ../../HW/src/dp/dp_fetch.vhd:953:61  */
  assign n7853_o = n7852_o & n7849_o;
  /* ../../HW/src/dp/dp_fetch.vhd:951:42  */
  assign n7854_o = n7853_o & bus_write_in;
  /* ../../HW/src/dp/dp_fetch.vhd:951:20  */
  assign n7855_o = n7854_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:959:44  */
  assign n7860_o = wregno == 5'b01000;
  /* ../../HW/src/dp/dp_fetch.vhd:959:34  */
  assign n7861_o = n7860_o & bus_write_r;
  /* ../../HW/src/dp/dp_fetch.vhd:959:81  */
  assign n7863_o = wregno2_r == 6'b010011;
  /* ../../HW/src/dp/dp_fetch.vhd:959:68  */
  assign n7864_o = n7863_o & n7861_o;
  /* ../../HW/src/dp/dp_fetch.vhd:959:13  */
  assign n7865_o = n7864_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:980:69  */
  assign n7869_o = print_param_rr[63:32];
  /* ../../HW/src/dp/dp_fetch.vhd:982:72  */
  assign n7871_o = print_param_rr[29:0];
  /* ../../HW/src/dp/dp_fetch.vhd:985:65  */
  assign n7872_o = task_busy_in[0];
  /* ../../HW/src/dp/dp_fetch.vhd:986:65  */
  assign n7873_o = task_busy_in[1];
  /* ../../HW/src/dp/dp_fetch.vhd:987:85  */
  assign n7874_o = sink_pcore_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:988:86  */
  assign n7875_o = pcore_source_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:989:80  */
  assign n7876_o = sink_sram_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:990:81  */
  assign n7877_o = sram_source_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:991:85  */
  assign n7878_o = sink_pcore_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:992:86  */
  assign n7879_o = pcore_source_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:993:80  */
  assign n7880_o = sink_sram_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:994:81  */
  assign n7881_o = sram_source_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:997:99  */
  assign n7882_o = log_time_r[19:0];
  assign n7885_o = n7883_o[31:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1009:19  */
  assign n7886_o = log_write[43:32];
  /* ../../HW/src/dp/dp_fetch.vhd:1009:93  */
  assign n7887_o = log_status_last_r[43:32];
  /* ../../HW/src/dp/dp_fetch.vhd:1009:73  */
  assign n7888_o = n7886_o != n7887_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1009:7  */
  assign n7891_o = n7888_o ? 1'b1 : 1'b0;
  assign n7892_o = {n7885_o, 2'b11};
  /* ../../HW/src/dp/dp_fetch.vhd:1002:4  */
  assign n7893_o = log2_valid_in ? log2_in : n7892_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1002:4  */
  assign n7895_o = log2_valid_in ? 1'b1 : n7891_o;
  /* ../../HW/src/dp/dp_fetch.vhd:998:4  */
  assign n7896_o = log1_valid_in ? log1_in : n7893_o;
  /* ../../HW/src/dp/dp_fetch.vhd:998:4  */
  assign n7898_o = log1_valid_in ? 1'b1 : n7895_o;
  assign n7899_o = {n7882_o, ddr_source_busy_r, sink_ddr_busy_r, n7881_o, n7880_o, n7879_o, n7878_o, n7877_o, n7876_o, n7875_o, n7874_o, n7873_o, n7872_o, n7896_o};
  assign n7900_o = {n7869_o, n7871_o, 2'b10};
  /* ../../HW/src/dp/dp_fetch.vhd:977:1  */
  assign n7901_o = print_indication_rr ? n7900_o : n7899_o;
  /* ../../HW/src/dp/dp_fetch.vhd:977:1  */
  assign n7903_o = print_indication_rr ? 1'b1 : n7898_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1024:25  */
  assign n7905_o = log_wrreq & log_enable_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1024:47  */
  assign n7906_o = ~log_full;
  /* ../../HW/src/dp/dp_fetch.vhd:1024:42  */
  assign n7907_o = n7905_o & n7906_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1040:14  */
  assign log_fifo_i_n7908 = log_fifo_i_q_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1043:18  */
  assign log_fifo_i_n7911 = log_fifo_i_empty_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1044:17  */
  assign log_fifo_i_n7912 = log_fifo_i_full_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1026:1  */
  scfifo_64_8_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 log_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(log_write),
    .write_in(log_wrreq2),
    .read_in(log_rdreq),
    .q_out(log_fifo_i_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(log_fifo_i_empty_out),
    .full_out(log_fifo_i_full_out),
    .almost_full_out());
  /* ../../HW/src/dp/dp_fetch.vhd:1056:56  */
  assign n7924_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1056:47  */
  assign n7925_o = n7924_o & ready;
  /* ../../HW/src/dp/dp_fetch.vhd:1056:31  */
  assign n7926_o = n7925_o & valid;
  /* ../../HW/src/dp/dp_fetch.vhd:1056:14  */
  assign n7927_o = n7926_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1064:24  */
  assign fifo_i_n7929 = fifo_i_readdata1_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1065:24  */
  assign fifo_i_n7930 = fifo_i_readdata2_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1066:26  */
  assign n7931_o = rdreqs[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1067:26  */
  assign n7932_o = rdreqs[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1068:21  */
  assign fifo_i_n7933 = fifo_i_valid1_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1069:21  */
  assign fifo_i_n7934 = fifo_i_valid2_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1070:19  */
  assign fifo_i_n7935 = fifo_i_full_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1071:27  */
  assign fifo_i_n7936 = fifo_i_fifo_avail_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1058:1  */
  dp_fifo fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .writedata_in(data),
    .wreq_in(wreq),
    .rdreq1_in(n7931_o),
    .rdreq2_in(n7932_o),
    .readdata1_out(fifo_i_readdata1_out),
    .readdata2_out(fifo_i_readdata2_out),
    .valid1_out(fifo_i_valid1_out),
    .valid2_out(fifo_i_valid2_out),
    .full_out(fifo_i_full_out),
    .fifo_avail_out(fifo_i_fifo_avail_out));
  /* ../../HW/src/dp/dp_fetch.vhd:1093:14  */
  assign gen1_ram_i_n7949 = gen1_ram_i_q_b; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1079:1  */
  ramw2_16_16_4_4_776_776 gen1_ram_i (
    .clock(clock_in),
    .clock_x2(clock_x2_in),
    .address_a(dp_var_waddress),
    .data_a(dp_var_write),
    .wren_a(dp_var_we),
    .address_b(dp_var_raddress),
    .q_b(gen1_ram_i_q_b));
  /* ../../HW/src/dp/dp_fetch.vhd:261:101  */
  assign n7959_o = template_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:263:107  */
  assign n7962_o = template_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:265:105  */
  assign n7964_o = template_r[72:48];
  /* ../../HW/src/dp/dp_fetch.vhd:267:105  */
  assign n7966_o = template_r[97:73];
  /* ../../HW/src/dp/dp_fetch.vhd:269:101  */
  assign n7968_o = template_r[121:98];
  /* ../../HW/src/dp/dp_fetch.vhd:271:107  */
  assign n7970_o = template_r[145:122];
  /* ../../HW/src/dp/dp_fetch.vhd:273:105  */
  assign n7972_o = template_r[170:146];
  /* ../../HW/src/dp/dp_fetch.vhd:275:105  */
  assign n7974_o = template_r[195:171];
  /* ../../HW/src/dp/dp_fetch.vhd:277:101  */
  assign n7976_o = template_r[219:196];
  /* ../../HW/src/dp/dp_fetch.vhd:279:107  */
  assign n7978_o = template_r[243:220];
  /* ../../HW/src/dp/dp_fetch.vhd:281:105  */
  assign n7980_o = template_r[268:244];
  /* ../../HW/src/dp/dp_fetch.vhd:283:105  */
  assign n7982_o = template_r[293:269];
  /* ../../HW/src/dp/dp_fetch.vhd:285:101  */
  assign n7984_o = template_r[317:294];
  /* ../../HW/src/dp/dp_fetch.vhd:287:107  */
  assign n7986_o = template_r[341:318];
  /* ../../HW/src/dp/dp_fetch.vhd:289:105  */
  assign n7988_o = template_r[366:342];
  /* ../../HW/src/dp/dp_fetch.vhd:291:105  */
  assign n7990_o = template_r[391:367];
  /* ../../HW/src/dp/dp_fetch.vhd:293:101  */
  assign n7992_o = template_r[415:392];
  /* ../../HW/src/dp/dp_fetch.vhd:295:107  */
  assign n7994_o = template_r[439:416];
  /* ../../HW/src/dp/dp_fetch.vhd:297:105  */
  assign n7996_o = template_r[464:440];
  /* ../../HW/src/dp/dp_fetch.vhd:299:105  */
  assign n7998_o = template_r[489:465];
  /* ../../HW/src/dp/dp_fetch.vhd:301:103  */
  assign n8000_o = template_r[514:490];
  /* ../../HW/src/dp/dp_fetch.vhd:303:104  */
  assign n8002_o = template_r[539:515];
  /* ../../HW/src/dp/dp_fetch.vhd:305:108  */
  assign n8004_o = template_r[564:540];
  /* ../../HW/src/dp/dp_fetch.vhd:307:109  */
  assign n8006_o = template_r[567:565];
  /* ../../HW/src/dp/dp_fetch.vhd:309:103  */
  assign n8008_o = template_r[592:568];
  /* ../../HW/src/dp/dp_fetch.vhd:311:97  */
  assign n8010_o = template_r[624:593];
  /* ../../HW/src/dp/dp_fetch.vhd:313:99  */
  assign n8012_o = template_r[648:625];
  /* ../../HW/src/dp/dp_fetch.vhd:315:105  */
  assign n8014_o = template_r[672:649];
  /* ../../HW/src/dp/dp_fetch.vhd:317:38  */
  assign n8016_o = template_r[673];
  /* ../../HW/src/dp/dp_fetch.vhd:319:104  */
  assign n8018_o = template_r[675:674];
  /* ../../HW/src/dp/dp_fetch.vhd:321:38  */
  assign n8020_o = template_r[676];
  /* ../../HW/src/dp/dp_fetch.vhd:323:104  */
  assign n8022_o = template_r[700:677];
  /* ../../HW/src/dp/dp_fetch.vhd:325:99  */
  assign n8024_o = template_r[706:701];
  /* ../../HW/src/dp/dp_fetch.vhd:327:98  */
  assign n8026_o = template_r[722:707];
  /* ../../HW/src/dp/dp_fetch.vhd:329:38  */
  assign n8028_o = template_r[723];
  /* ../../HW/src/dp/dp_fetch.vhd:331:102  */
  assign n8030_o = template_r[725:724];
  /* ../../HW/src/dp/dp_fetch.vhd:333:100  */
  assign n8032_o = template_r[727:726];
  /* ../../HW/src/dp/dp_fetch.vhd:335:101  */
  assign n8034_o = template_r[751:728];
  /* ../../HW/src/dp/dp_fetch.vhd:337:107  */
  assign n8036_o = template_r[775:752];
  assign n8037_o = {n7959_o, n7962_o, n7964_o, n7966_o, n7968_o, n7970_o, n7972_o, n7974_o, n7976_o, n7978_o, n7980_o, n7982_o, n7984_o, n7986_o, n7988_o, n7990_o, n7992_o, n7994_o, n7996_o, n7998_o, n8000_o, n8002_o, n8004_o, n8006_o, n8008_o, n8010_o, n8012_o, n8014_o, n8016_o, n8018_o, n8020_o, n8022_o, n8024_o, n8026_o, n8028_o, n8030_o, n8032_o, n8034_o, n8036_o};
  /* ../../HW/src/dp/dp_fetch.vhd:351:35  */
  assign n8045_o = dp_var_read[775:752];
  /* ../../HW/src/dp/dp_fetch.vhd:353:41  */
  assign n8048_o = dp_var_read[751:728];
  /* ../../HW/src/dp/dp_fetch.vhd:355:39  */
  assign n8050_o = dp_var_read[727:703];
  /* ../../HW/src/dp/dp_fetch.vhd:357:39  */
  assign n8052_o = dp_var_read[702:678];
  /* ../../HW/src/dp/dp_fetch.vhd:359:35  */
  assign n8054_o = dp_var_read[677:654];
  /* ../../HW/src/dp/dp_fetch.vhd:361:41  */
  assign n8056_o = dp_var_read[653:630];
  /* ../../HW/src/dp/dp_fetch.vhd:363:39  */
  assign n8058_o = dp_var_read[629:605];
  /* ../../HW/src/dp/dp_fetch.vhd:365:39  */
  assign n8060_o = dp_var_read[604:580];
  /* ../../HW/src/dp/dp_fetch.vhd:367:35  */
  assign n8062_o = dp_var_read[579:556];
  /* ../../HW/src/dp/dp_fetch.vhd:369:41  */
  assign n8064_o = dp_var_read[555:532];
  /* ../../HW/src/dp/dp_fetch.vhd:371:39  */
  assign n8066_o = dp_var_read[531:507];
  /* ../../HW/src/dp/dp_fetch.vhd:373:39  */
  assign n8068_o = dp_var_read[506:482];
  /* ../../HW/src/dp/dp_fetch.vhd:375:35  */
  assign n8070_o = dp_var_read[481:458];
  /* ../../HW/src/dp/dp_fetch.vhd:377:41  */
  assign n8072_o = dp_var_read[457:434];
  /* ../../HW/src/dp/dp_fetch.vhd:379:39  */
  assign n8074_o = dp_var_read[433:409];
  /* ../../HW/src/dp/dp_fetch.vhd:381:39  */
  assign n8076_o = dp_var_read[408:384];
  /* ../../HW/src/dp/dp_fetch.vhd:383:35  */
  assign n8078_o = dp_var_read[383:360];
  /* ../../HW/src/dp/dp_fetch.vhd:385:41  */
  assign n8080_o = dp_var_read[359:336];
  /* ../../HW/src/dp/dp_fetch.vhd:387:39  */
  assign n8082_o = dp_var_read[335:311];
  /* ../../HW/src/dp/dp_fetch.vhd:389:39  */
  assign n8084_o = dp_var_read[310:286];
  /* ../../HW/src/dp/dp_fetch.vhd:391:37  */
  assign n8086_o = dp_var_read[285:261];
  /* ../../HW/src/dp/dp_fetch.vhd:393:38  */
  assign n8088_o = dp_var_read[260:236];
  /* ../../HW/src/dp/dp_fetch.vhd:395:42  */
  assign n8090_o = dp_var_read[235:211];
  /* ../../HW/src/dp/dp_fetch.vhd:397:43  */
  assign n8092_o = dp_var_read[210:208];
  /* ../../HW/src/dp/dp_fetch.vhd:399:37  */
  assign n8094_o = dp_var_read[207:183];
  /* ../../HW/src/dp/dp_fetch.vhd:401:31  */
  assign n8096_o = dp_var_read[182:151];
  /* ../../HW/src/dp/dp_fetch.vhd:403:33  */
  assign n8098_o = dp_var_read[150:127];
  /* ../../HW/src/dp/dp_fetch.vhd:405:39  */
  assign n8100_o = dp_var_read[126:103];
  /* ../../HW/src/dp/dp_fetch.vhd:407:35  */
  assign n8102_o = dp_var_read[102];
  /* ../../HW/src/dp/dp_fetch.vhd:409:29  */
  assign n8104_o = dp_var_read[101:100];
  /* ../../HW/src/dp/dp_fetch.vhd:411:26  */
  assign n8106_o = dp_var_read[99];
  /* ../../HW/src/dp/dp_fetch.vhd:413:38  */
  assign n8108_o = dp_var_read[98:75];
  /* ../../HW/src/dp/dp_fetch.vhd:415:24  */
  assign n8110_o = dp_var_read[74:69];
  /* ../../HW/src/dp/dp_fetch.vhd:417:23  */
  assign n8112_o = dp_var_read[68:53];
  /* ../../HW/src/dp/dp_fetch.vhd:419:25  */
  assign n8114_o = dp_var_read[52];
  /* ../../HW/src/dp/dp_fetch.vhd:421:36  */
  assign n8116_o = dp_var_read[51:50];
  /* ../../HW/src/dp/dp_fetch.vhd:423:34  */
  assign n8118_o = dp_var_read[49:48];
  /* ../../HW/src/dp/dp_fetch.vhd:425:35  */
  assign n8120_o = dp_var_read[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:427:41  */
  assign n8122_o = dp_var_read[23:0];
  assign n8123_o = {n8122_o, n8120_o, n8118_o, n8116_o, n8114_o, n8112_o, n8110_o, n8108_o, n8106_o, n8104_o, n8102_o, n8100_o, n8098_o, n8096_o, n8094_o, n8092_o, n8090_o, n8088_o, n8086_o, n8084_o, n8082_o, n8080_o, n8078_o, n8076_o, n8074_o, n8072_o, n8070_o, n8068_o, n8066_o, n8064_o, n8062_o, n8060_o, n8058_o, n8056_o, n8054_o, n8052_o, n8050_o, n8048_o, n8045_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1123:44  */
  assign n8124_o = wregno2[3:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1123:95  */
  assign n8125_o = wregno2[3];
  /* ../../HW/src/dp/dp_fetch.vhd:1123:82  */
  assign n8126_o = n8125_o ? n8124_o : n8128_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1125:45  */
  assign n8127_o = wregno2[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1125:83  */
  assign n8128_o = {n8127_o, curr_vm_r};
  /* ../../HW/src/dp/dp_fetch.vhd:1131:48  */
  assign n8129_o = orec_generic[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1131:71  */
  assign n8130_o = orec_generic[96:33];
  /* ../../HW/src/dp/dp_fetch.vhd:1131:56  */
  assign n8131_o = {n8129_o, n8130_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1147:16  */
  assign indication_i_n8132 = indication_i_q_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1148:21  */
  assign indication_i_n8133 = indication_i_ravail_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1149:20  */
  assign indication_i_n8134 = indication_i_wused_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1150:20  */
  assign indication_i_n8135 = indication_i_empty_out; // (signal)
  /* ../../HW/src/dp/dp_fetch.vhd:1133:1  */
  scfifo_67_8_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 indication_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(in_indication),
    .write_in(wreq2_indication),
    .read_in(indication_rdreq),
    .q_out(indication_i_q_out),
    .ravail_out(indication_i_ravail_out),
    .wused_out(indication_i_wused_out),
    .empty_out(indication_i_empty_out),
    .full_out(),
    .almost_full_out());
  /* ../../HW/src/dp/dp_fetch.vhd:1156:48  */
  assign n8149_o = pcore_read_pending_p0_in | pcore_read_pending_p1_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1158:46  */
  assign n8150_o = sram_read_pending_p0_in | sram_read_pending_p1_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1160:44  */
  assign n8151_o = ddr_read_pending_p0_in | ddr_read_pending_p1_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1166:31  */
  assign n8152_o = bus_waddr_r[4:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1168:33  */
  assign n8153_o = bus_waddr_in[10:5];
  /* ../../HW/src/dp/dp_fetch.vhd:1170:34  */
  assign n8154_o = bus_waddr_r[10:5];
  /* ../../HW/src/dp/dp_fetch.vhd:1172:31  */
  assign n8155_o = bus_raddr_r[4:0];
  /* ../../HW/src/dp/dp_fetch.vhd:441:100  */
  assign n8166_o = irec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:443:103  */
  assign n8169_o = irec[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:445:38  */
  assign n8171_o = irec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:447:108  */
  assign n8173_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:447:115  */
  assign n8174_o = n8173_o[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:449:114  */
  assign n8176_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:449:121  */
  assign n8177_o = n8176_o[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:451:112  */
  assign n8179_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:451:119  */
  assign n8180_o = n8179_o[72:48];
  /* ../../HW/src/dp/dp_fetch.vhd:453:112  */
  assign n8182_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:453:119  */
  assign n8183_o = n8182_o[97:73];
  /* ../../HW/src/dp/dp_fetch.vhd:455:108  */
  assign n8185_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:455:115  */
  assign n8186_o = n8185_o[121:98];
  /* ../../HW/src/dp/dp_fetch.vhd:457:114  */
  assign n8188_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:457:121  */
  assign n8189_o = n8188_o[145:122];
  /* ../../HW/src/dp/dp_fetch.vhd:459:112  */
  assign n8191_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:459:119  */
  assign n8192_o = n8191_o[170:146];
  /* ../../HW/src/dp/dp_fetch.vhd:461:112  */
  assign n8194_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:461:119  */
  assign n8195_o = n8194_o[195:171];
  /* ../../HW/src/dp/dp_fetch.vhd:463:108  */
  assign n8197_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:463:115  */
  assign n8198_o = n8197_o[219:196];
  /* ../../HW/src/dp/dp_fetch.vhd:465:114  */
  assign n8200_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:465:121  */
  assign n8201_o = n8200_o[243:220];
  /* ../../HW/src/dp/dp_fetch.vhd:467:112  */
  assign n8203_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:467:119  */
  assign n8204_o = n8203_o[268:244];
  /* ../../HW/src/dp/dp_fetch.vhd:469:112  */
  assign n8206_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:469:119  */
  assign n8207_o = n8206_o[293:269];
  /* ../../HW/src/dp/dp_fetch.vhd:471:108  */
  assign n8209_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:471:115  */
  assign n8210_o = n8209_o[317:294];
  /* ../../HW/src/dp/dp_fetch.vhd:473:114  */
  assign n8212_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:473:121  */
  assign n8213_o = n8212_o[341:318];
  /* ../../HW/src/dp/dp_fetch.vhd:475:112  */
  assign n8215_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:475:119  */
  assign n8216_o = n8215_o[366:342];
  /* ../../HW/src/dp/dp_fetch.vhd:477:112  */
  assign n8218_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:477:119  */
  assign n8219_o = n8218_o[391:367];
  /* ../../HW/src/dp/dp_fetch.vhd:479:108  */
  assign n8221_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:479:115  */
  assign n8222_o = n8221_o[415:392];
  /* ../../HW/src/dp/dp_fetch.vhd:481:114  */
  assign n8224_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:481:121  */
  assign n8225_o = n8224_o[439:416];
  /* ../../HW/src/dp/dp_fetch.vhd:483:112  */
  assign n8227_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:483:119  */
  assign n8228_o = n8227_o[464:440];
  /* ../../HW/src/dp/dp_fetch.vhd:485:112  */
  assign n8230_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:485:119  */
  assign n8231_o = n8230_o[489:465];
  /* ../../HW/src/dp/dp_fetch.vhd:487:110  */
  assign n8233_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:487:117  */
  assign n8234_o = n8233_o[514:490];
  /* ../../HW/src/dp/dp_fetch.vhd:489:111  */
  assign n8236_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:489:118  */
  assign n8237_o = n8236_o[539:515];
  /* ../../HW/src/dp/dp_fetch.vhd:491:115  */
  assign n8239_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:491:122  */
  assign n8240_o = n8239_o[564:540];
  /* ../../HW/src/dp/dp_fetch.vhd:493:116  */
  assign n8242_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:493:123  */
  assign n8243_o = n8242_o[567:565];
  /* ../../HW/src/dp/dp_fetch.vhd:495:110  */
  assign n8245_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:495:117  */
  assign n8246_o = n8245_o[592:568];
  /* ../../HW/src/dp/dp_fetch.vhd:497:38  */
  assign n8248_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:497:45  */
  assign n8249_o = n8248_o[673];
  /* ../../HW/src/dp/dp_fetch.vhd:499:111  */
  assign n8251_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:499:118  */
  assign n8252_o = n8251_o[675:674];
  /* ../../HW/src/dp/dp_fetch.vhd:501:38  */
  assign n8254_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:501:45  */
  assign n8255_o = n8254_o[676];
  /* ../../HW/src/dp/dp_fetch.vhd:503:104  */
  assign n8257_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:503:111  */
  assign n8258_o = n8257_o[624:593];
  /* ../../HW/src/dp/dp_fetch.vhd:505:106  */
  assign n8260_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:505:113  */
  assign n8261_o = n8260_o[648:625];
  /* ../../HW/src/dp/dp_fetch.vhd:507:112  */
  assign n8263_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:507:119  */
  assign n8264_o = n8263_o[672:649];
  /* ../../HW/src/dp/dp_fetch.vhd:509:108  */
  assign n8266_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:509:115  */
  assign n8267_o = n8266_o[751:728];
  /* ../../HW/src/dp/dp_fetch.vhd:511:114  */
  assign n8269_o = irec[783:8];
  /* ../../HW/src/dp/dp_fetch.vhd:511:121  */
  assign n8270_o = n8269_o[775:752];
  /* ../../HW/src/dp/dp_fetch.vhd:513:107  */
  assign n8272_o = irec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:515:110  */
  assign n8274_o = irec[787:786];
  /* ../../HW/src/dp/dp_fetch.vhd:517:106  */
  assign n8276_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:517:111  */
  assign n8277_o = n8276_o[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:519:112  */
  assign n8279_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:519:117  */
  assign n8280_o = n8279_o[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:521:110  */
  assign n8282_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:521:115  */
  assign n8283_o = n8282_o[72:48];
  /* ../../HW/src/dp/dp_fetch.vhd:523:110  */
  assign n8285_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:523:115  */
  assign n8286_o = n8285_o[97:73];
  /* ../../HW/src/dp/dp_fetch.vhd:525:106  */
  assign n8288_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:525:111  */
  assign n8289_o = n8288_o[121:98];
  /* ../../HW/src/dp/dp_fetch.vhd:527:112  */
  assign n8291_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:527:117  */
  assign n8292_o = n8291_o[145:122];
  /* ../../HW/src/dp/dp_fetch.vhd:529:110  */
  assign n8294_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:529:115  */
  assign n8295_o = n8294_o[170:146];
  /* ../../HW/src/dp/dp_fetch.vhd:531:110  */
  assign n8297_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:531:115  */
  assign n8298_o = n8297_o[195:171];
  /* ../../HW/src/dp/dp_fetch.vhd:533:106  */
  assign n8300_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:533:111  */
  assign n8301_o = n8300_o[219:196];
  /* ../../HW/src/dp/dp_fetch.vhd:535:112  */
  assign n8303_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:535:117  */
  assign n8304_o = n8303_o[243:220];
  /* ../../HW/src/dp/dp_fetch.vhd:537:110  */
  assign n8306_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:537:115  */
  assign n8307_o = n8306_o[268:244];
  /* ../../HW/src/dp/dp_fetch.vhd:539:110  */
  assign n8309_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:539:115  */
  assign n8310_o = n8309_o[293:269];
  /* ../../HW/src/dp/dp_fetch.vhd:541:106  */
  assign n8312_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:541:111  */
  assign n8313_o = n8312_o[317:294];
  /* ../../HW/src/dp/dp_fetch.vhd:543:112  */
  assign n8315_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:543:117  */
  assign n8316_o = n8315_o[341:318];
  /* ../../HW/src/dp/dp_fetch.vhd:545:110  */
  assign n8318_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:545:115  */
  assign n8319_o = n8318_o[366:342];
  /* ../../HW/src/dp/dp_fetch.vhd:547:110  */
  assign n8321_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:547:115  */
  assign n8322_o = n8321_o[391:367];
  /* ../../HW/src/dp/dp_fetch.vhd:549:106  */
  assign n8324_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:549:111  */
  assign n8325_o = n8324_o[415:392];
  /* ../../HW/src/dp/dp_fetch.vhd:551:112  */
  assign n8327_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:551:117  */
  assign n8328_o = n8327_o[439:416];
  /* ../../HW/src/dp/dp_fetch.vhd:553:110  */
  assign n8330_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:553:115  */
  assign n8331_o = n8330_o[464:440];
  /* ../../HW/src/dp/dp_fetch.vhd:555:110  */
  assign n8333_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:555:115  */
  assign n8334_o = n8333_o[489:465];
  /* ../../HW/src/dp/dp_fetch.vhd:557:108  */
  assign n8336_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:557:113  */
  assign n8337_o = n8336_o[514:490];
  /* ../../HW/src/dp/dp_fetch.vhd:559:109  */
  assign n8339_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:559:114  */
  assign n8340_o = n8339_o[539:515];
  /* ../../HW/src/dp/dp_fetch.vhd:561:113  */
  assign n8342_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:561:118  */
  assign n8343_o = n8342_o[564:540];
  /* ../../HW/src/dp/dp_fetch.vhd:563:114  */
  assign n8345_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:563:119  */
  assign n8346_o = n8345_o[567:565];
  /* ../../HW/src/dp/dp_fetch.vhd:565:108  */
  assign n8348_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:565:113  */
  assign n8349_o = n8348_o[592:568];
  /* ../../HW/src/dp/dp_fetch.vhd:567:38  */
  assign n8351_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:567:43  */
  assign n8352_o = n8351_o[673];
  /* ../../HW/src/dp/dp_fetch.vhd:569:109  */
  assign n8354_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:569:114  */
  assign n8355_o = n8354_o[675:674];
  /* ../../HW/src/dp/dp_fetch.vhd:571:38  */
  assign n8357_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:571:43  */
  assign n8358_o = n8357_o[676];
  /* ../../HW/src/dp/dp_fetch.vhd:573:102  */
  assign n8360_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:573:107  */
  assign n8361_o = n8360_o[624:593];
  /* ../../HW/src/dp/dp_fetch.vhd:575:104  */
  assign n8363_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:575:109  */
  assign n8364_o = n8363_o[648:625];
  /* ../../HW/src/dp/dp_fetch.vhd:577:110  */
  assign n8366_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:577:115  */
  assign n8367_o = n8366_o[672:649];
  /* ../../HW/src/dp/dp_fetch.vhd:579:106  */
  assign n8369_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:579:111  */
  assign n8370_o = n8369_o[751:728];
  /* ../../HW/src/dp/dp_fetch.vhd:581:112  */
  assign n8372_o = irec[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:581:117  */
  assign n8373_o = n8372_o[775:752];
  /* ../../HW/src/dp/dp_fetch.vhd:583:105  */
  assign n8375_o = irec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:585:108  */
  assign n8377_o = irec[1567:1566];
  /* ../../HW/src/dp/dp_fetch.vhd:587:99  */
  assign n8379_o = irec[1573:1568];
  /* ../../HW/src/dp/dp_fetch.vhd:589:99  */
  assign n8381_o = irec[1597:1574];
  /* ../../HW/src/dp/dp_fetch.vhd:591:98  */
  assign n8383_o = irec[1613:1598];
  /* ../../HW/src/dp/dp_fetch.vhd:593:48  */
  assign n8385_o = irec[1614];
  /* ../../HW/src/dp/dp_fetch.vhd:595:48  */
  assign n8387_o = irec[1615];
  /* ../../HW/src/dp/dp_fetch.vhd:597:48  */
  assign n8389_o = irec[1616];
  /* ../../HW/src/dp/dp_fetch.vhd:599:48  */
  assign n8391_o = irec[1617];
  /* ../../HW/src/dp/dp_fetch.vhd:601:98  */
  assign n8393_o = irec[1619:1618];
  assign n8394_o = {n8166_o, n8169_o, n8171_o, n8174_o, n8177_o, n8180_o, n8183_o, n8186_o, n8189_o, n8192_o, n8195_o, n8198_o, n8201_o, n8204_o, n8207_o, n8210_o, n8213_o, n8216_o, n8219_o, n8222_o, n8225_o, n8228_o, n8231_o, n8234_o, n8237_o, n8240_o, n8243_o, n8246_o, n8249_o, n8252_o, n8255_o, n8258_o, n8261_o, n8264_o, n8267_o, n8270_o, n8272_o, n8274_o, n8277_o, n8280_o, n8283_o, n8286_o, n8289_o, n8292_o, n8295_o, n8298_o, n8301_o, n8304_o, n8307_o, n8310_o, n8313_o, n8316_o, n8319_o, n8322_o, n8325_o, n8328_o, n8331_o, n8334_o, n8337_o, n8340_o, n8343_o, n8346_o, n8349_o, n8352_o, n8355_o, n8358_o, n8361_o, n8364_o, n8367_o, n8370_o, n8373_o, n8375_o, n8377_o, n8379_o, n8381_o, n8383_o, n8385_o, n8387_o, n8389_o, n8391_o, n8393_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1182:36  */
  assign n8395_o = irec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1182:42  */
  assign n8397_o = n8395_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1182:25  */
  assign n8398_o = n8397_o ? n8394_o : n8416_o;
  /* ../../HW/src/dp/dp_fetch.vhd:789:35  */
  assign n8406_o = irec_generic[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:790:35  */
  assign n8407_o = irec_generic[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:789:43  */
  assign n8408_o = {n8406_o, n8407_o};
  /* ../../HW/src/dp/dp_fetch.vhd:791:18  */
  assign n8409_o = irec_generic[7];
  /* ../../HW/src/dp/dp_fetch.vhd:790:46  */
  assign n8410_o = {n8408_o, n8409_o};
  /* ../../HW/src/dp/dp_fetch.vhd:792:35  */
  assign n8411_o = irec_generic[32:8];
  /* ../../HW/src/dp/dp_fetch.vhd:791:21  */
  assign n8412_o = {n8410_o, n8411_o};
  /* ../../HW/src/dp/dp_fetch.vhd:793:35  */
  assign n8413_o = irec_generic[96:33];
  /* ../../HW/src/dp/dp_fetch.vhd:792:42  */
  assign n8414_o = {n8412_o, n8413_o};
  /* ../../HW/src/dp/dp_fetch.vhd:793:47  */
  assign n8416_o = {n8414_o, 1421'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
  /* ../../HW/src/dp/dp_fetch.vhd:615:34  */
  assign n8425_o = q1[1517:1515];
  /* ../../HW/src/dp/dp_fetch.vhd:617:28  */
  assign n8428_o = q1[1514:1511];
  /* ../../HW/src/dp/dp_fetch.vhd:619:21  */
  assign n8430_o = q1[1510];
  /* ../../HW/src/dp/dp_fetch.vhd:621:42  */
  assign n8432_o = q1[1509:1486];
  /* ../../HW/src/dp/dp_fetch.vhd:623:48  */
  assign n8434_o = q1[1485:1462];
  /* ../../HW/src/dp/dp_fetch.vhd:625:46  */
  assign n8436_o = q1[1461:1437];
  /* ../../HW/src/dp/dp_fetch.vhd:627:46  */
  assign n8438_o = q1[1436:1412];
  /* ../../HW/src/dp/dp_fetch.vhd:629:42  */
  assign n8440_o = q1[1411:1388];
  /* ../../HW/src/dp/dp_fetch.vhd:631:48  */
  assign n8442_o = q1[1387:1364];
  /* ../../HW/src/dp/dp_fetch.vhd:633:46  */
  assign n8444_o = q1[1363:1339];
  /* ../../HW/src/dp/dp_fetch.vhd:635:46  */
  assign n8446_o = q1[1338:1314];
  /* ../../HW/src/dp/dp_fetch.vhd:637:42  */
  assign n8448_o = q1[1313:1290];
  /* ../../HW/src/dp/dp_fetch.vhd:639:48  */
  assign n8450_o = q1[1289:1266];
  /* ../../HW/src/dp/dp_fetch.vhd:641:46  */
  assign n8452_o = q1[1265:1241];
  /* ../../HW/src/dp/dp_fetch.vhd:643:46  */
  assign n8454_o = q1[1240:1216];
  /* ../../HW/src/dp/dp_fetch.vhd:645:42  */
  assign n8456_o = q1[1215:1192];
  /* ../../HW/src/dp/dp_fetch.vhd:647:48  */
  assign n8458_o = q1[1191:1168];
  /* ../../HW/src/dp/dp_fetch.vhd:649:46  */
  assign n8460_o = q1[1167:1143];
  /* ../../HW/src/dp/dp_fetch.vhd:651:46  */
  assign n8462_o = q1[1142:1118];
  /* ../../HW/src/dp/dp_fetch.vhd:653:42  */
  assign n8464_o = q1[1117:1094];
  /* ../../HW/src/dp/dp_fetch.vhd:655:48  */
  assign n8466_o = q1[1093:1070];
  /* ../../HW/src/dp/dp_fetch.vhd:657:46  */
  assign n8468_o = q1[1069:1045];
  /* ../../HW/src/dp/dp_fetch.vhd:659:46  */
  assign n8470_o = q1[1044:1020];
  /* ../../HW/src/dp/dp_fetch.vhd:661:44  */
  assign n8472_o = q1[1019:995];
  /* ../../HW/src/dp/dp_fetch.vhd:663:45  */
  assign n8474_o = q1[994:970];
  /* ../../HW/src/dp/dp_fetch.vhd:665:49  */
  assign n8476_o = q1[969:945];
  /* ../../HW/src/dp/dp_fetch.vhd:667:50  */
  assign n8478_o = q1[944:942];
  /* ../../HW/src/dp/dp_fetch.vhd:669:44  */
  assign n8480_o = q1[941:917];
  /* ../../HW/src/dp/dp_fetch.vhd:671:42  */
  assign n8482_o = q1[916];
  /* ../../HW/src/dp/dp_fetch.vhd:673:36  */
  assign n8485_o = q1[915:914];
  /* ../../HW/src/dp/dp_fetch.vhd:675:33  */
  assign n8487_o = q1[913];
  /* ../../HW/src/dp/dp_fetch.vhd:677:38  */
  assign n8489_o = q1[912:881];
  /* ../../HW/src/dp/dp_fetch.vhd:679:40  */
  assign n8491_o = q1[880:857];
  /* ../../HW/src/dp/dp_fetch.vhd:681:46  */
  assign n8493_o = q1[856:833];
  /* ../../HW/src/dp/dp_fetch.vhd:683:42  */
  assign n8494_o = q1[832:809];
  assign n8496_o = n8426_o[735:685];
  /* ../../HW/src/dp/dp_fetch.vhd:685:48  */
  assign n8497_o = q1[808:785];
  /* ../../HW/src/dp/dp_fetch.vhd:687:41  */
  assign n8499_o = q1[784:783];
  /* ../../HW/src/dp/dp_fetch.vhd:689:44  */
  assign n8501_o = q1[782:781];
  /* ../../HW/src/dp/dp_fetch.vhd:691:40  */
  assign n8503_o = q1[780:757];
  /* ../../HW/src/dp/dp_fetch.vhd:693:46  */
  assign n8505_o = q1[756:733];
  /* ../../HW/src/dp/dp_fetch.vhd:695:44  */
  assign n8507_o = q1[732:708];
  /* ../../HW/src/dp/dp_fetch.vhd:697:44  */
  assign n8509_o = q1[707:683];
  /* ../../HW/src/dp/dp_fetch.vhd:699:40  */
  assign n8511_o = q1[682:659];
  /* ../../HW/src/dp/dp_fetch.vhd:701:46  */
  assign n8513_o = q1[658:635];
  /* ../../HW/src/dp/dp_fetch.vhd:703:44  */
  assign n8515_o = q1[634:610];
  /* ../../HW/src/dp/dp_fetch.vhd:705:44  */
  assign n8517_o = q1[609:585];
  /* ../../HW/src/dp/dp_fetch.vhd:707:40  */
  assign n8519_o = q1[584:561];
  /* ../../HW/src/dp/dp_fetch.vhd:709:46  */
  assign n8521_o = q1[560:537];
  /* ../../HW/src/dp/dp_fetch.vhd:711:44  */
  assign n8523_o = q1[536:512];
  /* ../../HW/src/dp/dp_fetch.vhd:713:44  */
  assign n8525_o = q1[511:487];
  /* ../../HW/src/dp/dp_fetch.vhd:715:40  */
  assign n8527_o = q1[486:463];
  /* ../../HW/src/dp/dp_fetch.vhd:717:46  */
  assign n8529_o = q1[462:439];
  /* ../../HW/src/dp/dp_fetch.vhd:719:44  */
  assign n8531_o = q1[438:414];
  /* ../../HW/src/dp/dp_fetch.vhd:721:44  */
  assign n8533_o = q1[413:389];
  /* ../../HW/src/dp/dp_fetch.vhd:723:40  */
  assign n8535_o = q1[388:365];
  /* ../../HW/src/dp/dp_fetch.vhd:725:46  */
  assign n8537_o = q1[364:341];
  /* ../../HW/src/dp/dp_fetch.vhd:727:44  */
  assign n8539_o = q1[340:316];
  /* ../../HW/src/dp/dp_fetch.vhd:729:44  */
  assign n8541_o = q1[315:291];
  /* ../../HW/src/dp/dp_fetch.vhd:731:42  */
  assign n8543_o = q1[290:266];
  /* ../../HW/src/dp/dp_fetch.vhd:733:43  */
  assign n8545_o = q1[265:241];
  /* ../../HW/src/dp/dp_fetch.vhd:735:47  */
  assign n8547_o = q1[240:216];
  /* ../../HW/src/dp/dp_fetch.vhd:737:48  */
  assign n8549_o = q1[215:213];
  /* ../../HW/src/dp/dp_fetch.vhd:739:42  */
  assign n8551_o = q1[212:188];
  /* ../../HW/src/dp/dp_fetch.vhd:741:40  */
  assign n8553_o = q1[187];
  /* ../../HW/src/dp/dp_fetch.vhd:743:34  */
  assign n8556_o = q1[186:185];
  /* ../../HW/src/dp/dp_fetch.vhd:745:31  */
  assign n8558_o = q1[184];
  /* ../../HW/src/dp/dp_fetch.vhd:747:36  */
  assign n8560_o = q1[183:152];
  /* ../../HW/src/dp/dp_fetch.vhd:749:38  */
  assign n8562_o = q1[151:128];
  /* ../../HW/src/dp/dp_fetch.vhd:751:44  */
  assign n8564_o = q1[127:104];
  /* ../../HW/src/dp/dp_fetch.vhd:753:40  */
  assign n8565_o = q1[103:80];
  assign n8567_o = n8426_o[1515:1465];
  /* ../../HW/src/dp/dp_fetch.vhd:755:46  */
  assign n8568_o = q1[79:56];
  /* ../../HW/src/dp/dp_fetch.vhd:757:39  */
  assign n8570_o = q1[55:54];
  /* ../../HW/src/dp/dp_fetch.vhd:759:42  */
  assign n8572_o = q1[53:52];
  /* ../../HW/src/dp/dp_fetch.vhd:761:24  */
  assign n8574_o = q1[51:46];
  /* ../../HW/src/dp/dp_fetch.vhd:763:33  */
  assign n8576_o = q1[45:22];
  /* ../../HW/src/dp/dp_fetch.vhd:765:23  */
  assign n8578_o = q1[21:6];
  /* ../../HW/src/dp/dp_fetch.vhd:767:25  */
  assign n8580_o = q1[5];
  /* ../../HW/src/dp/dp_fetch.vhd:769:35  */
  assign n8582_o = q1[4];
  /* ../../HW/src/dp/dp_fetch.vhd:771:33  */
  assign n8584_o = q1[3];
  /* ../../HW/src/dp/dp_fetch.vhd:773:33  */
  assign n8586_o = q1[2];
  /* ../../HW/src/dp/dp_fetch.vhd:775:45  */
  assign n8588_o = q1[1:0];
  assign n8589_o = {n8588_o, n8586_o, n8584_o, n8582_o, n8580_o, n8578_o, n8576_o, n8574_o, n8572_o, n8570_o, n8568_o, n8565_o, n8567_o, n8558_o, n8556_o, n8553_o, n8564_o, n8562_o, n8560_o, n8551_o, n8549_o, n8547_o, n8545_o, n8543_o, n8541_o, n8539_o, n8537_o, n8535_o, n8533_o, n8531_o, n8529_o, n8527_o, n8525_o, n8523_o, n8521_o, n8519_o, n8517_o, n8515_o, n8513_o, n8511_o, n8509_o, n8507_o, n8505_o, n8503_o, n8501_o, n8499_o, n8497_o, n8494_o, n8496_o, n8487_o, n8485_o, n8482_o, n8493_o, n8491_o, n8489_o, n8480_o, n8478_o, n8476_o, n8474_o, n8472_o, n8470_o, n8468_o, n8466_o, n8464_o, n8462_o, n8460_o, n8458_o, n8456_o, n8454_o, n8452_o, n8450_o, n8448_o, n8446_o, n8444_o, n8442_o, n8440_o, n8438_o, n8436_o, n8434_o, n8432_o, n8430_o, n8428_o, n8425_o};
  /* ../../HW/src/dp/dp_fetch.vhd:615:34  */
  assign n8597_o = q2[1517:1515];
  /* ../../HW/src/dp/dp_fetch.vhd:617:28  */
  assign n8600_o = q2[1514:1511];
  /* ../../HW/src/dp/dp_fetch.vhd:619:21  */
  assign n8602_o = q2[1510];
  /* ../../HW/src/dp/dp_fetch.vhd:621:42  */
  assign n8604_o = q2[1509:1486];
  /* ../../HW/src/dp/dp_fetch.vhd:623:48  */
  assign n8606_o = q2[1485:1462];
  /* ../../HW/src/dp/dp_fetch.vhd:625:46  */
  assign n8608_o = q2[1461:1437];
  /* ../../HW/src/dp/dp_fetch.vhd:627:46  */
  assign n8610_o = q2[1436:1412];
  /* ../../HW/src/dp/dp_fetch.vhd:629:42  */
  assign n8612_o = q2[1411:1388];
  /* ../../HW/src/dp/dp_fetch.vhd:631:48  */
  assign n8614_o = q2[1387:1364];
  /* ../../HW/src/dp/dp_fetch.vhd:633:46  */
  assign n8616_o = q2[1363:1339];
  /* ../../HW/src/dp/dp_fetch.vhd:635:46  */
  assign n8618_o = q2[1338:1314];
  /* ../../HW/src/dp/dp_fetch.vhd:637:42  */
  assign n8620_o = q2[1313:1290];
  /* ../../HW/src/dp/dp_fetch.vhd:639:48  */
  assign n8622_o = q2[1289:1266];
  /* ../../HW/src/dp/dp_fetch.vhd:641:46  */
  assign n8624_o = q2[1265:1241];
  /* ../../HW/src/dp/dp_fetch.vhd:643:46  */
  assign n8626_o = q2[1240:1216];
  /* ../../HW/src/dp/dp_fetch.vhd:645:42  */
  assign n8628_o = q2[1215:1192];
  /* ../../HW/src/dp/dp_fetch.vhd:647:48  */
  assign n8630_o = q2[1191:1168];
  /* ../../HW/src/dp/dp_fetch.vhd:649:46  */
  assign n8632_o = q2[1167:1143];
  /* ../../HW/src/dp/dp_fetch.vhd:651:46  */
  assign n8634_o = q2[1142:1118];
  /* ../../HW/src/dp/dp_fetch.vhd:653:42  */
  assign n8636_o = q2[1117:1094];
  /* ../../HW/src/dp/dp_fetch.vhd:655:48  */
  assign n8638_o = q2[1093:1070];
  /* ../../HW/src/dp/dp_fetch.vhd:657:46  */
  assign n8640_o = q2[1069:1045];
  /* ../../HW/src/dp/dp_fetch.vhd:659:46  */
  assign n8642_o = q2[1044:1020];
  /* ../../HW/src/dp/dp_fetch.vhd:661:44  */
  assign n8644_o = q2[1019:995];
  /* ../../HW/src/dp/dp_fetch.vhd:663:45  */
  assign n8646_o = q2[994:970];
  /* ../../HW/src/dp/dp_fetch.vhd:665:49  */
  assign n8648_o = q2[969:945];
  /* ../../HW/src/dp/dp_fetch.vhd:667:50  */
  assign n8650_o = q2[944:942];
  /* ../../HW/src/dp/dp_fetch.vhd:669:44  */
  assign n8652_o = q2[941:917];
  /* ../../HW/src/dp/dp_fetch.vhd:671:42  */
  assign n8654_o = q2[916];
  /* ../../HW/src/dp/dp_fetch.vhd:673:36  */
  assign n8657_o = q2[915:914];
  /* ../../HW/src/dp/dp_fetch.vhd:675:33  */
  assign n8659_o = q2[913];
  /* ../../HW/src/dp/dp_fetch.vhd:677:38  */
  assign n8661_o = q2[912:881];
  /* ../../HW/src/dp/dp_fetch.vhd:679:40  */
  assign n8663_o = q2[880:857];
  /* ../../HW/src/dp/dp_fetch.vhd:681:46  */
  assign n8665_o = q2[856:833];
  /* ../../HW/src/dp/dp_fetch.vhd:683:42  */
  assign n8666_o = q2[832:809];
  assign n8668_o = n8598_o[735:685];
  /* ../../HW/src/dp/dp_fetch.vhd:685:48  */
  assign n8669_o = q2[808:785];
  /* ../../HW/src/dp/dp_fetch.vhd:687:41  */
  assign n8671_o = q2[784:783];
  /* ../../HW/src/dp/dp_fetch.vhd:689:44  */
  assign n8673_o = q2[782:781];
  /* ../../HW/src/dp/dp_fetch.vhd:691:40  */
  assign n8675_o = q2[780:757];
  /* ../../HW/src/dp/dp_fetch.vhd:693:46  */
  assign n8677_o = q2[756:733];
  /* ../../HW/src/dp/dp_fetch.vhd:695:44  */
  assign n8679_o = q2[732:708];
  /* ../../HW/src/dp/dp_fetch.vhd:697:44  */
  assign n8681_o = q2[707:683];
  /* ../../HW/src/dp/dp_fetch.vhd:699:40  */
  assign n8683_o = q2[682:659];
  /* ../../HW/src/dp/dp_fetch.vhd:701:46  */
  assign n8685_o = q2[658:635];
  /* ../../HW/src/dp/dp_fetch.vhd:703:44  */
  assign n8687_o = q2[634:610];
  /* ../../HW/src/dp/dp_fetch.vhd:705:44  */
  assign n8689_o = q2[609:585];
  /* ../../HW/src/dp/dp_fetch.vhd:707:40  */
  assign n8691_o = q2[584:561];
  /* ../../HW/src/dp/dp_fetch.vhd:709:46  */
  assign n8693_o = q2[560:537];
  /* ../../HW/src/dp/dp_fetch.vhd:711:44  */
  assign n8695_o = q2[536:512];
  /* ../../HW/src/dp/dp_fetch.vhd:713:44  */
  assign n8697_o = q2[511:487];
  /* ../../HW/src/dp/dp_fetch.vhd:715:40  */
  assign n8699_o = q2[486:463];
  /* ../../HW/src/dp/dp_fetch.vhd:717:46  */
  assign n8701_o = q2[462:439];
  /* ../../HW/src/dp/dp_fetch.vhd:719:44  */
  assign n8703_o = q2[438:414];
  /* ../../HW/src/dp/dp_fetch.vhd:721:44  */
  assign n8705_o = q2[413:389];
  /* ../../HW/src/dp/dp_fetch.vhd:723:40  */
  assign n8707_o = q2[388:365];
  /* ../../HW/src/dp/dp_fetch.vhd:725:46  */
  assign n8709_o = q2[364:341];
  /* ../../HW/src/dp/dp_fetch.vhd:727:44  */
  assign n8711_o = q2[340:316];
  /* ../../HW/src/dp/dp_fetch.vhd:729:44  */
  assign n8713_o = q2[315:291];
  /* ../../HW/src/dp/dp_fetch.vhd:731:42  */
  assign n8715_o = q2[290:266];
  /* ../../HW/src/dp/dp_fetch.vhd:733:43  */
  assign n8717_o = q2[265:241];
  /* ../../HW/src/dp/dp_fetch.vhd:735:47  */
  assign n8719_o = q2[240:216];
  /* ../../HW/src/dp/dp_fetch.vhd:737:48  */
  assign n8721_o = q2[215:213];
  /* ../../HW/src/dp/dp_fetch.vhd:739:42  */
  assign n8723_o = q2[212:188];
  /* ../../HW/src/dp/dp_fetch.vhd:741:40  */
  assign n8725_o = q2[187];
  /* ../../HW/src/dp/dp_fetch.vhd:743:34  */
  assign n8728_o = q2[186:185];
  /* ../../HW/src/dp/dp_fetch.vhd:745:31  */
  assign n8730_o = q2[184];
  /* ../../HW/src/dp/dp_fetch.vhd:747:36  */
  assign n8732_o = q2[183:152];
  /* ../../HW/src/dp/dp_fetch.vhd:749:38  */
  assign n8734_o = q2[151:128];
  /* ../../HW/src/dp/dp_fetch.vhd:751:44  */
  assign n8736_o = q2[127:104];
  /* ../../HW/src/dp/dp_fetch.vhd:753:40  */
  assign n8737_o = q2[103:80];
  assign n8739_o = n8598_o[1515:1465];
  /* ../../HW/src/dp/dp_fetch.vhd:755:46  */
  assign n8740_o = q2[79:56];
  /* ../../HW/src/dp/dp_fetch.vhd:757:39  */
  assign n8742_o = q2[55:54];
  /* ../../HW/src/dp/dp_fetch.vhd:759:42  */
  assign n8744_o = q2[53:52];
  /* ../../HW/src/dp/dp_fetch.vhd:761:24  */
  assign n8746_o = q2[51:46];
  /* ../../HW/src/dp/dp_fetch.vhd:763:33  */
  assign n8748_o = q2[45:22];
  /* ../../HW/src/dp/dp_fetch.vhd:765:23  */
  assign n8750_o = q2[21:6];
  /* ../../HW/src/dp/dp_fetch.vhd:767:25  */
  assign n8752_o = q2[5];
  /* ../../HW/src/dp/dp_fetch.vhd:769:35  */
  assign n8754_o = q2[4];
  /* ../../HW/src/dp/dp_fetch.vhd:771:33  */
  assign n8756_o = q2[3];
  /* ../../HW/src/dp/dp_fetch.vhd:773:33  */
  assign n8758_o = q2[2];
  /* ../../HW/src/dp/dp_fetch.vhd:775:45  */
  assign n8760_o = q2[1:0];
  assign n8761_o = {n8760_o, n8758_o, n8756_o, n8754_o, n8752_o, n8750_o, n8748_o, n8746_o, n8744_o, n8742_o, n8740_o, n8737_o, n8739_o, n8730_o, n8728_o, n8725_o, n8736_o, n8734_o, n8732_o, n8723_o, n8721_o, n8719_o, n8717_o, n8715_o, n8713_o, n8711_o, n8709_o, n8707_o, n8705_o, n8703_o, n8701_o, n8699_o, n8697_o, n8695_o, n8693_o, n8691_o, n8689_o, n8687_o, n8685_o, n8683_o, n8681_o, n8679_o, n8677_o, n8675_o, n8673_o, n8671_o, n8669_o, n8666_o, n8668_o, n8659_o, n8657_o, n8654_o, n8665_o, n8663_o, n8661_o, n8652_o, n8650_o, n8648_o, n8646_o, n8644_o, n8642_o, n8640_o, n8638_o, n8636_o, n8634_o, n8632_o, n8630_o, n8628_o, n8626_o, n8624_o, n8622_o, n8620_o, n8618_o, n8616_o, n8614_o, n8612_o, n8610_o, n8608_o, n8606_o, n8604_o, n8602_o, n8600_o, n8597_o};
  /* ../../HW/src/dp/dp_fetch.vhd:807:34  */
  assign n8769_o = q1[1517:1515];
  /* ../../HW/src/dp/dp_fetch.vhd:809:28  */
  assign n8772_o = q1[1514:1511];
  /* ../../HW/src/dp/dp_fetch.vhd:811:21  */
  assign n8774_o = q1[1510];
  /* ../../HW/src/dp/dp_fetch.vhd:813:24  */
  assign n8776_o = q1[1509:1485];
  /* ../../HW/src/dp/dp_fetch.vhd:815:29  */
  assign n8778_o = q1[1484:1421];
  assign n8779_o = {n8778_o, n8776_o, n8774_o, n8772_o, n8769_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1197:43  */
  assign n8781_o = src_template_r[725:724];
  /* ../../HW/src/dp/dp_fetch.vhd:1197:67  */
  assign n8782_o = src_template_r[727:726];
  /* ../../HW/src/dp/dp_fetch.vhd:1197:90  */
  assign n8783_o = dest_template_r[727:726];
  /* ../../HW/src/dp/dp_fetch.vhd:1198:44  */
  assign n8784_o = dest_template_r[706:701];
  /* ../../HW/src/dp/dp_fetch.vhd:1198:66  */
  assign n8785_o = dest_template_r[700:677];
  /* ../../HW/src/dp/dp_fetch.vhd:1199:43  */
  assign n8786_o = src_template_r[722:707];
  /* ../../HW/src/dp/dp_fetch.vhd:1199:63  */
  assign n8787_o = src_template_r[723];
  /* ../../HW/src/dp/dp_fetch.vhd:840:45  */
  assign n8795_o = bus_writedata_r[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:842:35  */
  assign n8798_o = bus_writedata_r[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:857:46  */
  assign n8808_o = bus_writedata_r[14];
  /* ../../HW/src/dp/dp_fetch.vhd:859:44  */
  assign n8811_o = bus_writedata_r[15];
  /* ../../HW/src/dp/dp_fetch.vhd:861:44  */
  assign n8813_o = bus_writedata_r[16];
  /* ../../HW/src/dp/dp_fetch.vhd:863:56  */
  assign n8815_o = bus_writedata_r[18:17];
  assign n8819_o = {n8815_o, n8813_o, n8811_o, n8808_o, n8787_o, n8786_o, n8785_o, n8784_o, n8781_o, n8783_o, dest_template_r, n8781_o, n8782_o, src_template_r, curr_vm_r, n8798_o, n8795_o};
  /* ../../HW/src/dp/dp_fetch.vhd:884:45  */
  assign n8827_o = bus_writedata_r[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:886:39  */
  assign n8830_o = bus_writedata_r[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:889:35  */
  assign n8833_o = bus_writedata_r[31:7];
  assign n8835_o = {indication_parm_r, n8833_o, curr_vm_r, n8830_o, n8827_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1208:33  */
  assign n8838_o = wregno == 5'b00101;
  /* ../../HW/src/dp/dp_fetch.vhd:1207:38  */
  assign n8839_o = n8838_o & bus_write_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1207:17  */
  assign n8840_o = n8839_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1212:19  */
  assign n8842_o = wreq_all & match;
  /* ../../HW/src/dp/dp_fetch.vhd:1221:42  */
  assign n8844_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1221:33  */
  assign n8845_o = n8844_o & valid;
  /* ../../HW/src/dp/dp_fetch.vhd:1221:60  */
  assign n8846_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1221:67  */
  assign n8848_o = n8846_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1221:50  */
  assign n8849_o = n8848_o & n8845_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1221:18  */
  assign n8850_o = n8849_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1223:42  */
  assign n8853_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1223:33  */
  assign n8854_o = n8853_o & valid;
  /* ../../HW/src/dp/dp_fetch.vhd:1223:60  */
  assign n8855_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1223:67  */
  assign n8857_o = n8855_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1223:50  */
  assign n8858_o = n8857_o & n8854_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1223:18  */
  assign n8859_o = n8858_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1227:27  */
  assign n8863_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1227:34  */
  assign n8865_o = n8863_o != 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1227:17  */
  assign n8866_o = n8865_o & valid;
  /* ../../HW/src/dp/dp_fetch.vhd:1230:16  */
  assign n8867_o = ready2[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1231:14  */
  assign n8868_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1231:46  */
  assign n8869_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1231:28  */
  assign n8870_o = n8868_o != n8869_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1231:59  */
  assign n8871_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1231:85  */
  assign n8872_o = dest_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1231:70  */
  assign n8873_o = n8871_o != n8872_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1231:50  */
  assign n8874_o = n8873_o & n8870_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1231:99  */
  assign n8875_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1231:90  */
  assign n8876_o = n8874_o | n8875_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1230:24  */
  assign n8877_o = n8876_o & n8867_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1233:22  */
  assign n8878_o = ready2[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1235:16  */
  assign n8879_o = ready2[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1236:17  */
  assign n8880_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1236:49  */
  assign n8881_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1236:31  */
  assign n8882_o = n8880_o != n8881_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1236:62  */
  assign n8883_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1236:88  */
  assign n8884_o = dest_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1236:73  */
  assign n8885_o = n8883_o != n8884_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1236:53  */
  assign n8886_o = n8885_o & n8882_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1236:102  */
  assign n8887_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1236:93  */
  assign n8888_o = n8886_o | n8887_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1235:24  */
  assign n8889_o = n8888_o & n8879_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1238:22  */
  assign n8890_o = ready2[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1235:4  */
  assign n8892_o = n8889_o ? n8890_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1235:4  */
  assign n8895_o = n8889_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1230:4  */
  assign n8896_o = n8877_o ? n8878_o : n8892_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1230:4  */
  assign n8898_o = n8877_o ? 1'b0 : n8895_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1227:4  */
  assign n8900_o = n8866_o ? 1'b1 : n8896_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1227:4  */
  assign n8902_o = n8866_o ? 1'b0 : n8898_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1246:55  */
  assign n8906_o = rregno == 5'b01011;
  /* ../../HW/src/dp/dp_fetch.vhd:1246:45  */
  assign n8907_o = n8906_o & bus_read_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1246:88  */
  assign n8908_o = match & n8907_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1246:25  */
  assign n8909_o = n8908_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1248:48  */
  assign n8913_o = rregno == 5'b00010;
  /* ../../HW/src/dp/dp_fetch.vhd:1248:38  */
  assign n8914_o = n8913_o & bus_read_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1248:74  */
  assign n8915_o = match & n8914_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1248:102  */
  assign n8916_o = ~log_empty;
  /* ../../HW/src/dp/dp_fetch.vhd:1248:88  */
  assign n8917_o = n8916_o & n8915_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1248:18  */
  assign n8918_o = n8917_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1256:15  */
  assign n8922_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1266:24  */
  assign n8924_o = ~waitrequest;
  /* ../../HW/src/dp/dp_fetch.vhd:1266:10  */
  assign n8926_o = n8924_o ? bus_write_in : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1285:17  */
  assign n8947_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1295:34  */
  assign n8950_o = indication[31:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1297:31  */
  assign n8951_o = match & bus_read_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1298:26  */
  assign n8953_o = rregno == 5'b01011;
  /* ../../HW/src/dp/dp_fetch.vhd:1301:47  */
  assign n8954_o = indication[63:32];
  /* ../../HW/src/dp/dp_fetch.vhd:1304:29  */
  assign n8956_o = rregno == 5'b01010;
  /* ../../HW/src/dp/dp_fetch.vhd:1308:29  */
  assign n8959_o = rregno == 5'b11001;
  /* ../../HW/src/dp/dp_fetch.vhd:1312:29  */
  assign n8961_o = rregno == 5'b01100;
  assign n8962_o = {24'b000000000000000000000000, indication_rdusedw};
  /* ../../HW/src/dp/dp_fetch.vhd:1316:29  */
  assign n8964_o = rregno == 5'b01110;
  /* ../../HW/src/dp/dp_fetch.vhd:1321:29  */
  assign n8967_o = rregno == 5'b00010;
  /* ../../HW/src/dp/dp_fetch.vhd:1322:33  */
  assign n8968_o = ~log_empty;
  /* ../../HW/src/dp/dp_fetch.vhd:1323:50  */
  assign n8969_o = log_read[31:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1322:21  */
  assign n8971_o = n8968_o ? n8969_o : 32'b00000000000000000000000000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:1327:47  */
  assign n8972_o = log_read[63:32];
  /* ../../HW/src/dp/dp_fetch.vhd:1329:29  */
  assign n8974_o = rregno == 5'b00011;
  /* ../../HW/src/dp/dp_fetch.vhd:1329:17  */
  assign n8976_o = n8974_o ? log_readtime_r : 32'b00000000000000000000000000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:1329:17  */
  assign n8979_o = n8974_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1321:17  */
  assign n8980_o = n8967_o ? n8971_o : n8976_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1321:17  */
  assign n8981_o = n8967_o ? n8972_o : log_readtime_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1321:17  */
  assign n8983_o = n8967_o ? 1'b1 : n8979_o;
  assign n8984_o = {24'b000000000000000000000000, fifo_avail};
  /* ../../HW/src/dp/dp_fetch.vhd:1316:17  */
  assign n8985_o = n8964_o ? n8984_o : n8980_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1316:17  */
  assign n8986_o = n8964_o ? log_readtime_r : n8981_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1316:17  */
  assign n8988_o = n8964_o ? 1'b1 : n8983_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1312:17  */
  assign n8989_o = n8961_o ? n8962_o : n8985_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1312:17  */
  assign n8990_o = n8961_o ? log_readtime_r : n8986_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1312:17  */
  assign n8992_o = n8961_o ? 1'b1 : n8988_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1308:17  */
  assign n8993_o = n8959_o ? indication_r : n8989_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1308:17  */
  assign n8994_o = n8959_o ? log_readtime_r : n8990_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1308:17  */
  assign n8996_o = n8959_o ? 1'b1 : n8992_o;
  assign n8997_o = {31'b0000000000000000000000000000000, indication_sync_r};
  /* ../../HW/src/dp/dp_fetch.vhd:1304:17  */
  assign n8998_o = n8956_o ? n8997_o : n8993_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1304:17  */
  assign n8999_o = n8956_o ? log_readtime_r : n8994_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1304:17  */
  assign n9001_o = n8956_o ? 1'b1 : n8996_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1298:17  */
  assign n9005_o = n8953_o ? n8950_o : n8998_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1298:17  */
  assign n9006_o = n8953_o ? log_readtime_r : n8999_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1298:17  */
  assign n9008_o = n8953_o ? 1'b1 : n9001_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1297:13  */
  assign n9009_o = n8953_o & n8951_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1297:13  */
  assign n9010_o = n8953_o & n8951_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1297:13  */
  assign n9014_o = n8951_o ? n9008_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1352:17  */
  assign n9046_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1364:32  */
  assign n9049_o = load_busid_r == 4'b1110;
  /* ../../HW/src/dp/dp_fetch.vhd:1366:35  */
  assign n9051_o = load_busid_r == 4'b1111;
  /* ../../HW/src/dp/dp_fetch.vhd:1366:17  */
  assign n9052_o = n9051_o ? template_r : dest_template_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1364:17  */
  assign n9054_o = n9049_o ? dest_template_r : n9052_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9055_o = n9049_o & load_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9058_o = load_r ? 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 : template_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1372:26  */
  assign n9060_o = wregno == 5'b01000;
  /* ../../HW/src/dp/dp_fetch.vhd:1374:33  */
  assign n9062_o = wregno2_r == 6'b000000;
  /* ../../HW/src/dp/dp_fetch.vhd:1375:71  */
  assign n9063_o = bus_writedata_r[23:0];
  assign n9064_o = n9057_o[23:0];
  assign n9065_o = template_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9066_o = load_r ? n9064_o : n9065_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1374:21  */
  assign n9067_o = n9062_o ? n9063_o : n9066_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1377:33  */
  assign n9069_o = wregno2_r == 6'b000001;
  /* ../../HW/src/dp/dp_fetch.vhd:1378:77  */
  assign n9070_o = bus_writedata_r[23:0];
  assign n9071_o = n9057_o[47:24];
  assign n9072_o = template_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9073_o = load_r ? n9071_o : n9072_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1377:21  */
  assign n9074_o = n9069_o ? n9070_o : n9073_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1380:33  */
  assign n9076_o = wregno2_r == 6'b001001;
  /* ../../HW/src/dp/dp_fetch.vhd:1381:75  */
  assign n9077_o = bus_writedata_r[24:0];
  assign n9078_o = n9057_o[72:48];
  assign n9079_o = template_r[72:48];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9080_o = load_r ? n9078_o : n9079_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1380:21  */
  assign n9081_o = n9076_o ? n9077_o : n9080_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1383:33  */
  assign n9083_o = wregno2_r == 6'b000010;
  /* ../../HW/src/dp/dp_fetch.vhd:1384:71  */
  assign n9084_o = bus_writedata_r[23:0];
  assign n9085_o = n9057_o[121:98];
  assign n9086_o = template_r[121:98];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9087_o = load_r ? n9085_o : n9086_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1383:21  */
  assign n9088_o = n9083_o ? n9084_o : n9087_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1386:33  */
  assign n9090_o = wregno2_r == 6'b000011;
  /* ../../HW/src/dp/dp_fetch.vhd:1387:77  */
  assign n9091_o = bus_writedata_r[23:0];
  assign n9092_o = n9057_o[145:122];
  assign n9093_o = template_r[145:122];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9094_o = load_r ? n9092_o : n9093_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1386:21  */
  assign n9095_o = n9090_o ? n9091_o : n9094_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1389:33  */
  assign n9097_o = wregno2_r == 6'b001010;
  /* ../../HW/src/dp/dp_fetch.vhd:1390:75  */
  assign n9098_o = bus_writedata_r[24:0];
  assign n9099_o = n9057_o[170:146];
  assign n9100_o = template_r[170:146];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9101_o = load_r ? n9099_o : n9100_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1389:21  */
  assign n9102_o = n9097_o ? n9098_o : n9101_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1392:33  */
  assign n9104_o = wregno2_r == 6'b000110;
  /* ../../HW/src/dp/dp_fetch.vhd:1393:71  */
  assign n9105_o = bus_writedata_r[23:0];
  assign n9106_o = n9057_o[219:196];
  assign n9107_o = template_r[219:196];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9108_o = load_r ? n9106_o : n9107_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1392:21  */
  assign n9109_o = n9104_o ? n9105_o : n9108_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1395:33  */
  assign n9111_o = wregno2_r == 6'b000111;
  /* ../../HW/src/dp/dp_fetch.vhd:1396:77  */
  assign n9112_o = bus_writedata_r[23:0];
  assign n9113_o = n9057_o[243:220];
  assign n9114_o = template_r[243:220];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9115_o = load_r ? n9113_o : n9114_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1395:21  */
  assign n9116_o = n9111_o ? n9112_o : n9115_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1398:33  */
  assign n9118_o = wregno2_r == 6'b001011;
  /* ../../HW/src/dp/dp_fetch.vhd:1399:75  */
  assign n9119_o = bus_writedata_r[24:0];
  assign n9120_o = n9057_o[268:244];
  assign n9121_o = template_r[268:244];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9122_o = load_r ? n9120_o : n9121_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1398:21  */
  assign n9123_o = n9118_o ? n9119_o : n9122_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1401:33  */
  assign n9125_o = wregno2_r == 6'b001101;
  /* ../../HW/src/dp/dp_fetch.vhd:1402:71  */
  assign n9126_o = bus_writedata_r[23:0];
  assign n9127_o = n9057_o[317:294];
  assign n9128_o = template_r[317:294];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9129_o = load_r ? n9127_o : n9128_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1401:21  */
  assign n9130_o = n9125_o ? n9126_o : n9129_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1404:33  */
  assign n9132_o = wregno2_r == 6'b001110;
  /* ../../HW/src/dp/dp_fetch.vhd:1405:77  */
  assign n9133_o = bus_writedata_r[23:0];
  assign n9134_o = n9057_o[341:318];
  assign n9135_o = template_r[341:318];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9136_o = load_r ? n9134_o : n9135_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1404:21  */
  assign n9137_o = n9132_o ? n9133_o : n9136_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1407:33  */
  assign n9139_o = wregno2_r == 6'b001111;
  /* ../../HW/src/dp/dp_fetch.vhd:1408:75  */
  assign n9140_o = bus_writedata_r[24:0];
  assign n9141_o = n9057_o[366:342];
  assign n9142_o = template_r[366:342];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9143_o = load_r ? n9141_o : n9142_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1407:21  */
  assign n9144_o = n9139_o ? n9140_o : n9143_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1410:33  */
  assign n9146_o = wregno2_r == 6'b010000;
  /* ../../HW/src/dp/dp_fetch.vhd:1411:71  */
  assign n9147_o = bus_writedata_r[23:0];
  assign n9148_o = n9057_o[415:392];
  assign n9149_o = template_r[415:392];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9150_o = load_r ? n9148_o : n9149_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1410:21  */
  assign n9151_o = n9146_o ? n9147_o : n9150_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1413:33  */
  assign n9153_o = wregno2_r == 6'b010001;
  /* ../../HW/src/dp/dp_fetch.vhd:1414:77  */
  assign n9154_o = bus_writedata_r[23:0];
  assign n9155_o = n9057_o[439:416];
  assign n9156_o = template_r[439:416];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9157_o = load_r ? n9155_o : n9156_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1413:21  */
  assign n9158_o = n9153_o ? n9154_o : n9157_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1416:33  */
  assign n9160_o = wregno2_r == 6'b010010;
  /* ../../HW/src/dp/dp_fetch.vhd:1417:75  */
  assign n9161_o = bus_writedata_r[24:0];
  assign n9162_o = n9057_o[464:440];
  assign n9163_o = template_r[464:440];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9164_o = load_r ? n9162_o : n9163_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1416:21  */
  assign n9165_o = n9160_o ? n9161_o : n9164_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1419:33  */
  assign n9167_o = wregno2_r == 6'b001100;
  /* ../../HW/src/dp/dp_fetch.vhd:1420:73  */
  assign n9168_o = bus_writedata_r[24:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1421:74  */
  assign n9169_o = bus_writedata_r[24:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1422:78  */
  assign n9170_o = bus_writedata_r[24:0];
  assign n9171_o = {n9170_o, n9169_o, n9168_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1424:33  */
  assign n9177_o = wregno2_r == 6'b011011;
  /* ../../HW/src/dp/dp_fetch.vhd:1425:74  */
  assign n9178_o = bus_writedata_r[24:0];
  assign n9179_o = n9171_o[49:25];
  assign n9180_o = n9057_o[539:515];
  assign n9181_o = template_r[539:515];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9182_o = load_r ? n9180_o : n9181_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1419:21  */
  assign n9183_o = n9167_o ? n9179_o : n9182_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1424:21  */
  assign n9184_o = n9177_o ? n9178_o : n9183_o;
  assign n9185_o = n9171_o[74:50];
  assign n9186_o = n9057_o[564:540];
  assign n9187_o = template_r[564:540];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9188_o = load_r ? n9186_o : n9187_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1419:21  */
  assign n9189_o = n9167_o ? n9185_o : n9188_o;
  assign n9190_o = n9171_o[24:0];
  assign n9191_o = n9057_o[514:490];
  assign n9192_o = template_r[514:490];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9193_o = load_r ? n9191_o : n9192_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1419:21  */
  assign n9194_o = n9167_o ? n9190_o : n9193_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1427:33  */
  assign n9196_o = wregno2_r == 6'b100000;
  /* ../../HW/src/dp/dp_fetch.vhd:1428:78  */
  assign n9197_o = bus_writedata_r[24:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1427:21  */
  assign n9198_o = n9196_o ? n9197_o : n9189_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1430:33  */
  assign n9200_o = wregno2_r == 6'b100001;
  /* ../../HW/src/dp/dp_fetch.vhd:1431:79  */
  assign n9201_o = bus_writedata_r[2:0];
  assign n9202_o = n9057_o[567:565];
  assign n9203_o = template_r[567:565];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9204_o = load_r ? n9202_o : n9203_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1430:21  */
  assign n9205_o = n9200_o ? n9201_o : n9204_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:33  */
  assign n9207_o = wregno2_r == 6'b000100;
  /* ../../HW/src/dp/dp_fetch.vhd:1437:58  */
  assign n9208_o = template_r[624:593];
  /* ../../HW/src/dp/dp_fetch.vhd:1437:61  */
  assign n9209_o = n9208_o + bus_writedata_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1440:33  */
  assign n9216_o = wregno2_r == 6'b011111;
  /* ../../HW/src/dp/dp_fetch.vhd:1441:71  */
  assign n9217_o = bus_writedata_r[23:0];
  assign n9218_o = n9057_o[751:728];
  assign n9219_o = template_r[751:728];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9220_o = load_r ? n9218_o : n9219_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1440:21  */
  assign n9221_o = n9216_o ? n9217_o : n9220_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1443:33  */
  assign n9223_o = wregno2_r == 6'b100010;
  /* ../../HW/src/dp/dp_fetch.vhd:1444:77  */
  assign n9224_o = bus_writedata_r[23:0];
  assign n9225_o = n9057_o[775:752];
  assign n9226_o = template_r[775:752];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9227_o = load_r ? n9225_o : n9226_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1443:21  */
  assign n9228_o = n9223_o ? n9224_o : n9227_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1446:33  */
  assign n9230_o = wregno2_r == 6'b000101;
  /* ../../HW/src/dp/dp_fetch.vhd:1447:69  */
  assign n9231_o = bus_writedata_r[23:0];
  assign n9232_o = n9057_o[648:625];
  assign n9233_o = template_r[648:625];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9234_o = load_r ? n9232_o : n9233_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1446:21  */
  assign n9235_o = n9230_o ? n9231_o : n9234_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1449:33  */
  assign n9237_o = wregno2_r == 6'b001000;
  /* ../../HW/src/dp/dp_fetch.vhd:1450:75  */
  assign n9238_o = bus_writedata_r[23:0];
  assign n9239_o = n9057_o[672:649];
  assign n9240_o = template_r[672:649];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9241_o = load_r ? n9239_o : n9240_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1449:21  */
  assign n9242_o = n9237_o ? n9238_o : n9241_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1452:33  */
  assign n9244_o = wregno2_r == 6'b010011;
  /* ../../HW/src/dp/dp_fetch.vhd:1453:43  */
  assign n9245_o = bus_writedata_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1455:74  */
  assign n9246_o = bus_writedata_r[5];
  /* ../../HW/src/dp/dp_fetch.vhd:1457:75  */
  assign n9247_o = bus_writedata_r[7:6];
  /* ../../HW/src/dp/dp_fetch.vhd:1459:68  */
  assign n9248_o = bus_writedata_r[9:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1461:65  */
  assign n9249_o = bus_writedata_r[10];
  /* ../../HW/src/dp/dp_fetch.vhd:1463:64  */
  assign n9250_o = bus_writedata_r[12:11];
  /* ../../HW/src/dp/dp_fetch.vhd:1465:39  */
  assign n9252_o = n9250_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:1467:42  */
  assign n9254_o = n9250_o == 2'b00;
  assign n9255_o = bus_writedata_r[21];
  assign n9256_o = n9209_o[21];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9257_o = load_r ? n9255_o : n9256_o;
  assign n9258_o = n9057_o[614];
  assign n9259_o = template_r[614];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9260_o = load_r ? n9258_o : n9259_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9261_o = n9207_o ? n9257_o : n9260_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1467:28  */
  assign n9262_o = n9254_o ? curr_vm_r : n9261_o;
  assign n9263_o = bus_writedata_r[14];
  assign n9264_o = n9209_o[14];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9265_o = load_r ? n9263_o : n9264_o;
  assign n9266_o = n9057_o[607];
  assign n9267_o = template_r[607];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9268_o = load_r ? n9266_o : n9267_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9269_o = n9207_o ? n9265_o : n9268_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1465:28  */
  assign n9270_o = n9252_o ? curr_vm_r : n9269_o;
  assign n9271_o = bus_writedata_r[21];
  assign n9272_o = n9209_o[21];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9273_o = load_r ? n9271_o : n9272_o;
  assign n9274_o = n9057_o[614];
  assign n9275_o = template_r[614];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9276_o = load_r ? n9274_o : n9275_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9277_o = n9207_o ? n9273_o : n9276_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1465:28  */
  assign n9278_o = n9252_o ? n9277_o : n9262_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1471:64  */
  assign n9279_o = bus_writedata_r[13];
  /* ../../HW/src/dp/dp_fetch.vhd:1473:63  */
  assign n9280_o = bus_writedata_r[19:14];
  assign n9281_o = {n9249_o, n9248_o, n9246_o};
  assign n9282_o = {n9250_o, n9247_o, n9279_o};
  assign n9283_o = bus_writedata_r[14];
  assign n9284_o = n9209_o[14];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9285_o = load_r ? n9283_o : n9284_o;
  assign n9286_o = n9057_o[607];
  assign n9287_o = template_r[607];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9288_o = load_r ? n9286_o : n9287_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9289_o = n9207_o ? n9285_o : n9288_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1453:25  */
  assign n9290_o = n9245_o ? n9270_o : n9289_o;
  assign n9291_o = bus_writedata_r[21];
  assign n9292_o = n9209_o[21];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9293_o = load_r ? n9291_o : n9292_o;
  assign n9294_o = n9057_o[614];
  assign n9295_o = template_r[614];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9296_o = load_r ? n9294_o : n9295_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9297_o = n9207_o ? n9293_o : n9296_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1453:25  */
  assign n9298_o = n9245_o ? n9278_o : n9297_o;
  assign n9299_o = n9057_o[676:673];
  assign n9300_o = template_r[676:673];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9301_o = load_r ? n9299_o : n9300_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1453:25  */
  assign n9302_o = n9245_o ? n9281_o : n9301_o;
  assign n9303_o = n9057_o[706:701];
  assign n9304_o = template_r[706:701];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9305_o = load_r ? n9303_o : n9304_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1453:25  */
  assign n9306_o = n9245_o ? n9280_o : n9305_o;
  assign n9307_o = n9057_o[727:723];
  assign n9308_o = template_r[727:723];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9309_o = load_r ? n9307_o : n9308_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1453:25  */
  assign n9310_o = n9245_o ? n9282_o : n9309_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1476:44  */
  assign n9314_o = bus_writedata_r[4];
  /* ../../HW/src/dp/dp_fetch.vhd:1477:68  */
  assign n9315_o = bus_writedata_r[4:1];
  /* ../../HW/src/dp/dp_fetch.vhd:1479:104  */
  assign n9316_o = bus_writedata_r[3:1];
  assign n9317_o = {n9316_o, curr_vm_r};
  /* ../../HW/src/dp/dp_fetch.vhd:1476:25  */
  assign n9318_o = n9314_o ? n9315_o : n9317_o;
  assign n9320_o = bus_writedata_r[14];
  assign n9321_o = n9209_o[14];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9322_o = load_r ? n9320_o : n9321_o;
  assign n9323_o = n9057_o[607];
  assign n9324_o = template_r[607];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9325_o = load_r ? n9323_o : n9324_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9326_o = n9207_o ? n9322_o : n9325_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1452:21  */
  assign n9327_o = n9244_o ? n9290_o : n9326_o;
  assign n9328_o = bus_writedata_r[21];
  assign n9329_o = n9209_o[21];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9330_o = load_r ? n9328_o : n9329_o;
  assign n9331_o = n9057_o[614];
  assign n9332_o = template_r[614];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9333_o = load_r ? n9331_o : n9332_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9334_o = n9207_o ? n9330_o : n9333_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1452:21  */
  assign n9335_o = n9244_o ? n9298_o : n9334_o;
  assign n9336_o = n9057_o[676:673];
  assign n9337_o = template_r[676:673];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9338_o = load_r ? n9336_o : n9337_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1452:21  */
  assign n9339_o = n9244_o ? n9302_o : n9338_o;
  assign n9340_o = n9057_o[706:701];
  assign n9341_o = template_r[706:701];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9342_o = load_r ? n9340_o : n9341_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1452:21  */
  assign n9343_o = n9244_o ? n9306_o : n9342_o;
  assign n9344_o = n9057_o[727:723];
  assign n9345_o = template_r[727:723];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9346_o = load_r ? n9344_o : n9345_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1452:21  */
  assign n9347_o = n9244_o ? n9310_o : n9346_o;
  assign n9355_o = bus_writedata_r[13:0];
  assign n9356_o = n9209_o[13:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9357_o = load_r ? n9355_o : n9356_o;
  assign n9358_o = n9057_o[606:593];
  assign n9359_o = template_r[606:593];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9360_o = load_r ? n9358_o : n9359_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9361_o = n9207_o ? n9357_o : n9360_o;
  assign n9362_o = bus_writedata_r[31:22];
  assign n9363_o = n9209_o[31:22];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9364_o = load_r ? n9362_o : n9363_o;
  assign n9365_o = n9057_o[624:615];
  assign n9366_o = template_r[624:615];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9367_o = load_r ? n9365_o : n9366_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9368_o = n9207_o ? n9364_o : n9367_o;
  assign n9369_o = bus_writedata_r[20:15];
  assign n9370_o = n9209_o[20:15];
  /* ../../HW/src/dp/dp_fetch.vhd:1434:25  */
  assign n9371_o = load_r ? n9369_o : n9370_o;
  assign n9372_o = n9057_o[613:608];
  assign n9373_o = template_r[613:608];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9374_o = load_r ? n9372_o : n9373_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1433:21  */
  assign n9375_o = n9207_o ? n9371_o : n9374_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1483:33  */
  assign n9379_o = wregno2_r == 6'b010100;
  /* ../../HW/src/dp/dp_fetch.vhd:1484:75  */
  assign n9380_o = bus_writedata_r[24:0];
  assign n9381_o = n9057_o[97:73];
  assign n9382_o = template_r[97:73];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9383_o = load_r ? n9381_o : n9382_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1483:21  */
  assign n9384_o = n9379_o ? n9380_o : n9383_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1486:33  */
  assign n9386_o = wregno2_r == 6'b010101;
  /* ../../HW/src/dp/dp_fetch.vhd:1487:75  */
  assign n9387_o = bus_writedata_r[24:0];
  assign n9388_o = n9057_o[195:171];
  assign n9389_o = template_r[195:171];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9390_o = load_r ? n9388_o : n9389_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1486:21  */
  assign n9391_o = n9386_o ? n9387_o : n9390_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1489:33  */
  assign n9393_o = wregno2_r == 6'b010110;
  /* ../../HW/src/dp/dp_fetch.vhd:1490:75  */
  assign n9394_o = bus_writedata_r[24:0];
  assign n9395_o = n9057_o[293:269];
  assign n9396_o = template_r[293:269];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9397_o = load_r ? n9395_o : n9396_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1489:21  */
  assign n9398_o = n9393_o ? n9394_o : n9397_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1492:33  */
  assign n9400_o = wregno2_r == 6'b010111;
  /* ../../HW/src/dp/dp_fetch.vhd:1493:75  */
  assign n9401_o = bus_writedata_r[24:0];
  assign n9402_o = n9057_o[391:367];
  assign n9403_o = template_r[391:367];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9404_o = load_r ? n9402_o : n9403_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1492:21  */
  assign n9405_o = n9400_o ? n9401_o : n9404_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1495:33  */
  assign n9407_o = wregno2_r == 6'b011000;
  /* ../../HW/src/dp/dp_fetch.vhd:1496:75  */
  assign n9408_o = bus_writedata_r[24:0];
  assign n9409_o = n9057_o[489:465];
  assign n9410_o = template_r[489:465];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9411_o = load_r ? n9409_o : n9410_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1495:21  */
  assign n9412_o = n9407_o ? n9408_o : n9411_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1498:33  */
  assign n9414_o = wregno2_r == 6'b011001;
  /* ../../HW/src/dp/dp_fetch.vhd:1499:73  */
  assign n9415_o = bus_writedata_r[24:0];
  assign n9416_o = n9057_o[592:568];
  assign n9417_o = template_r[592:568];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9418_o = load_r ? n9416_o : n9417_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1498:21  */
  assign n9419_o = n9414_o ? n9415_o : n9418_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1501:33  */
  assign n9421_o = wregno2_r == 6'b011010;
  /* ../../HW/src/dp/dp_fetch.vhd:1503:74  */
  assign n9422_o = bus_writedata_r[23:0];
  assign n9423_o = n9057_o[700:677];
  assign n9424_o = template_r[700:677];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9425_o = load_r ? n9423_o : n9424_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1501:21  */
  assign n9426_o = n9421_o ? n9422_o : n9425_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1505:33  */
  assign n9428_o = wregno2_r == 6'b011100;
  /* ../../HW/src/dp/dp_fetch.vhd:1507:59  */
  assign n9429_o = bus_writedata_r[15:0];
  assign n9430_o = n9057_o[722:707];
  assign n9431_o = template_r[722:707];
  /* ../../HW/src/dp/dp_fetch.vhd:1362:13  */
  assign n9432_o = load_r ? n9430_o : n9431_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1505:21  */
  assign n9433_o = n9428_o ? n9429_o : n9432_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1509:29  */
  assign n9435_o = wregno == 5'b01101;
  /* ../../HW/src/dp/dp_fetch.vhd:1509:17  */
  assign n9436_o = n9435_o ? dp_var_template : n9058_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1372:17  */
  assign n9437_o = n9244_o & n9060_o;
  assign n9438_o = {n9228_o, n9221_o, n9347_o, n9433_o, n9343_o, n9426_o, n9339_o, n9242_o, n9235_o, n9368_o, n9335_o, n9375_o, n9327_o, n9361_o, n9419_o, n9205_o, n9198_o, n9184_o, n9194_o, n9412_o, n9165_o, n9158_o, n9151_o, n9405_o, n9144_o, n9137_o, n9130_o, n9398_o, n9123_o, n9116_o, n9109_o, n9391_o, n9102_o, n9095_o, n9088_o, n9384_o, n9081_o, n9074_o, n9067_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1372:17  */
  assign n9439_o = n9060_o ? n9438_o : n9436_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1512:26  */
  assign n9443_o = wregno == 5'b10111;
  assign n9444_o = indication_parm_r[31:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1512:17  */
  assign n9445_o = n9443_o ? bus_writedata_r : n9444_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1516:26  */
  assign n9447_o = wregno == 5'b11000;
  assign n9448_o = indication_parm_r[63:32];
  /* ../../HW/src/dp/dp_fetch.vhd:1516:17  */
  assign n9449_o = n9447_o ? bus_writedata_r : n9448_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1520:26  */
  assign n9451_o = wregno == 5'b01001;
  /* ../../HW/src/dp/dp_fetch.vhd:1521:34  */
  assign n9452_o = ~curr_vm_r;
  assign n9454_o = {n9449_o, n9445_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1371:13  */
  assign n9456_o = n9437_o & bus_write_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1371:13  */
  assign n9457_o = n9451_o & bus_write_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1371:13  */
  assign n9458_o = bus_write_r ? n9439_o : n9058_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1524:13  */
  assign n9463_o = load ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1535:10  */
  always @*
    n9498_source_is_safe_v = n9766_o; // (isignal)
  initial
    n9498_source_is_safe_v = 16'bX;
  /* ../../HW/src/dp/dp_fetch.vhd:1536:10  */
  always @*
    n9498_dest_is_safe_v = n9785_o; // (isignal)
  initial
    n9498_dest_is_safe_v = 16'bX;
  /* ../../HW/src/dp/dp_fetch.vhd:1538:13  */
  assign n9502_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1547:93  */
  assign n9504_o = sram_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1547:72  */
  assign n9505_o = ~n9504_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1547:142  */
  assign n9506_o = ddr_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1547:122  */
  assign n9507_o = ~n9506_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1547:117  */
  assign n9508_o = n9505_o & n9507_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1548:90  */
  assign n9509_o = pcore_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1548:68  */
  assign n9510_o = ~n9509_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1548:139  */
  assign n9511_o = ddr_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1548:119  */
  assign n9512_o = ~n9511_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1548:114  */
  assign n9513_o = n9510_o & n9512_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1549:89  */
  assign n9514_o = pcore_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1549:67  */
  assign n9515_o = ~n9514_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1549:139  */
  assign n9516_o = sram_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1549:118  */
  assign n9517_o = ~n9516_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1549:113  */
  assign n9518_o = n9515_o & n9517_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1551:89  */
  assign n9519_o = sram_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1551:68  */
  assign n9520_o = ~n9519_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1551:134  */
  assign n9521_o = ddr_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1551:114  */
  assign n9522_o = ~n9521_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1551:109  */
  assign n9523_o = n9520_o & n9522_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1552:86  */
  assign n9524_o = pcore_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1552:64  */
  assign n9525_o = ~n9524_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1552:131  */
  assign n9526_o = ddr_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1552:111  */
  assign n9527_o = ~n9526_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1552:106  */
  assign n9528_o = n9525_o & n9527_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1553:85  */
  assign n9529_o = pcore_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1553:63  */
  assign n9530_o = ~n9529_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1553:131  */
  assign n9531_o = sram_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1553:110  */
  assign n9532_o = ~n9531_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1553:105  */
  assign n9533_o = n9530_o & n9532_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1555:88  */
  assign n9534_o = sram_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1555:67  */
  assign n9535_o = ~n9534_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1555:132  */
  assign n9536_o = ddr_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1555:112  */
  assign n9537_o = ~n9536_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1555:107  */
  assign n9538_o = n9535_o & n9537_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1556:85  */
  assign n9539_o = pcore_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1556:63  */
  assign n9540_o = ~n9539_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1556:129  */
  assign n9541_o = ddr_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1556:109  */
  assign n9542_o = ~n9541_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1556:104  */
  assign n9543_o = n9540_o & n9542_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1557:84  */
  assign n9544_o = pcore_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1557:62  */
  assign n9545_o = ~n9544_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1557:129  */
  assign n9546_o = sram_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1557:108  */
  assign n9547_o = ~n9546_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1557:103  */
  assign n9548_o = n9545_o & n9547_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1563:92  */
  assign n9549_o = pcore_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1563:70  */
  assign n9550_o = ~n9549_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1563:139  */
  assign n9551_o = pcore_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1563:117  */
  assign n9552_o = ~n9551_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1563:112  */
  assign n9553_o = n9550_o & n9552_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1564:88  */
  assign n9554_o = pcore_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1564:66  */
  assign n9555_o = ~n9554_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1564:139  */
  assign n9556_o = pcore_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1564:117  */
  assign n9557_o = ~n9556_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1564:112  */
  assign n9558_o = n9555_o & n9557_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1565:87  */
  assign n9559_o = pcore_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1565:65  */
  assign n9560_o = ~n9559_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1565:138  */
  assign n9561_o = pcore_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1565:116  */
  assign n9562_o = ~n9561_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1565:111  */
  assign n9563_o = n9560_o & n9562_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1567:87  */
  assign n9564_o = sram_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1567:66  */
  assign n9565_o = ~n9564_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1567:133  */
  assign n9566_o = sram_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1567:112  */
  assign n9567_o = ~n9566_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1567:107  */
  assign n9568_o = n9565_o & n9567_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1568:83  */
  assign n9569_o = sram_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1568:62  */
  assign n9570_o = ~n9569_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1568:133  */
  assign n9571_o = sram_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1568:112  */
  assign n9572_o = ~n9571_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1568:107  */
  assign n9573_o = n9570_o & n9572_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1569:82  */
  assign n9574_o = sram_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1569:61  */
  assign n9575_o = ~n9574_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1569:132  */
  assign n9576_o = sram_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1569:111  */
  assign n9577_o = ~n9576_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1569:106  */
  assign n9578_o = n9575_o & n9577_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1571:85  */
  assign n9579_o = ddr_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1571:65  */
  assign n9580_o = ~n9579_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1571:130  */
  assign n9581_o = ddr_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1571:110  */
  assign n9582_o = ~n9581_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1571:105  */
  assign n9583_o = n9580_o & n9582_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1572:81  */
  assign n9584_o = ddr_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1572:61  */
  assign n9585_o = ~n9584_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1572:130  */
  assign n9586_o = ddr_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1572:110  */
  assign n9587_o = ~n9586_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1572:105  */
  assign n9588_o = n9585_o & n9587_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1573:80  */
  assign n9589_o = ddr_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1573:60  */
  assign n9590_o = ~n9589_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1573:129  */
  assign n9591_o = ddr_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1573:109  */
  assign n9592_o = ~n9591_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1573:104  */
  assign n9593_o = n9590_o & n9592_o;
  assign n9594_o = n9498_source_is_safe_v[3];
  assign n9595_o = n9498_source_is_safe_v[7];
  assign n9596_o = n9498_source_is_safe_v[15:11];
  assign n9597_o = {n9596_o, n9548_o, n9543_o, n9538_o, n9595_o, n9533_o, n9528_o, n9523_o, n9594_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1576:110  */
  assign n9598_o = n9597_o[0];
  assign n9599_o = n9498_dest_is_safe_v[3];
  assign n9600_o = n9498_dest_is_safe_v[7];
  assign n9601_o = n9498_dest_is_safe_v[15:11];
  assign n9602_o = {n9601_o, n9593_o, n9588_o, n9583_o, n9600_o, n9578_o, n9573_o, n9568_o, n9599_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1576:173  */
  assign n9603_o = n9602_o[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1576:133  */
  assign n9604_o = n9598_o & n9603_o;
  assign n9605_o = n9498_source_is_safe_v[3];
  assign n9606_o = n9498_source_is_safe_v[7];
  assign n9607_o = n9498_source_is_safe_v[15:11];
  assign n9608_o = {n9607_o, n9548_o, n9543_o, n9538_o, n9606_o, n9533_o, n9528_o, n9523_o, n9605_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1577:106  */
  assign n9609_o = n9608_o[1];
  assign n9610_o = n9498_dest_is_safe_v[3];
  assign n9611_o = n9498_dest_is_safe_v[7];
  assign n9612_o = n9498_dest_is_safe_v[15:11];
  assign n9613_o = {n9612_o, n9593_o, n9588_o, n9583_o, n9611_o, n9578_o, n9573_o, n9568_o, n9610_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1577:161  */
  assign n9614_o = n9613_o[4];
  /* ../../HW/src/dp/dp_fetch.vhd:1577:125  */
  assign n9615_o = n9609_o & n9614_o;
  assign n9616_o = n9498_source_is_safe_v[3];
  assign n9617_o = n9498_source_is_safe_v[7];
  assign n9618_o = n9498_source_is_safe_v[15:11];
  assign n9619_o = {n9618_o, n9548_o, n9543_o, n9538_o, n9617_o, n9533_o, n9528_o, n9523_o, n9616_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1578:105  */
  assign n9620_o = n9619_o[2];
  assign n9621_o = n9498_dest_is_safe_v[3];
  assign n9622_o = n9498_dest_is_safe_v[7];
  assign n9623_o = n9498_dest_is_safe_v[15:11];
  assign n9624_o = {n9623_o, n9593_o, n9588_o, n9583_o, n9622_o, n9578_o, n9573_o, n9568_o, n9621_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1578:158  */
  assign n9625_o = n9624_o[8];
  /* ../../HW/src/dp/dp_fetch.vhd:1578:123  */
  assign n9626_o = n9620_o & n9625_o;
  assign n9627_o = n9498_source_is_safe_v[3];
  assign n9628_o = n9498_source_is_safe_v[7];
  assign n9629_o = n9498_source_is_safe_v[15:11];
  assign n9630_o = {n9629_o, n9548_o, n9543_o, n9538_o, n9628_o, n9533_o, n9528_o, n9523_o, n9627_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1579:102  */
  assign n9631_o = n9630_o[4];
  assign n9632_o = n9498_dest_is_safe_v[3];
  assign n9633_o = n9498_dest_is_safe_v[7];
  assign n9634_o = n9498_dest_is_safe_v[15:11];
  assign n9635_o = {n9634_o, n9593_o, n9588_o, n9583_o, n9633_o, n9578_o, n9573_o, n9568_o, n9632_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1579:165  */
  assign n9636_o = n9635_o[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1579:125  */
  assign n9637_o = n9631_o & n9636_o;
  assign n9638_o = n9498_source_is_safe_v[3];
  assign n9639_o = n9498_source_is_safe_v[7];
  assign n9640_o = n9498_source_is_safe_v[15:11];
  assign n9641_o = {n9640_o, n9548_o, n9543_o, n9538_o, n9639_o, n9533_o, n9528_o, n9523_o, n9638_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1580:98  */
  assign n9642_o = n9641_o[5];
  assign n9643_o = n9498_dest_is_safe_v[3];
  assign n9644_o = n9498_dest_is_safe_v[7];
  assign n9645_o = n9498_dest_is_safe_v[15:11];
  assign n9646_o = {n9645_o, n9593_o, n9588_o, n9583_o, n9644_o, n9578_o, n9573_o, n9568_o, n9643_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1580:153  */
  assign n9647_o = n9646_o[5];
  /* ../../HW/src/dp/dp_fetch.vhd:1580:117  */
  assign n9648_o = n9642_o & n9647_o;
  assign n9649_o = n9498_source_is_safe_v[3];
  assign n9650_o = n9498_source_is_safe_v[7];
  assign n9651_o = n9498_source_is_safe_v[15:11];
  assign n9652_o = {n9651_o, n9548_o, n9543_o, n9538_o, n9650_o, n9533_o, n9528_o, n9523_o, n9649_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1581:97  */
  assign n9653_o = n9652_o[6];
  assign n9654_o = n9498_dest_is_safe_v[3];
  assign n9655_o = n9498_dest_is_safe_v[7];
  assign n9656_o = n9498_dest_is_safe_v[15:11];
  assign n9657_o = {n9656_o, n9593_o, n9588_o, n9583_o, n9655_o, n9578_o, n9573_o, n9568_o, n9654_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1581:150  */
  assign n9658_o = n9657_o[9];
  /* ../../HW/src/dp/dp_fetch.vhd:1581:115  */
  assign n9659_o = n9653_o & n9658_o;
  assign n9660_o = n9498_source_is_safe_v[3];
  assign n9661_o = n9498_source_is_safe_v[7];
  assign n9662_o = n9498_source_is_safe_v[15:11];
  assign n9663_o = {n9662_o, n9548_o, n9543_o, n9538_o, n9661_o, n9533_o, n9528_o, n9523_o, n9660_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1582:100  */
  assign n9664_o = n9663_o[8];
  assign n9665_o = n9498_dest_is_safe_v[3];
  assign n9666_o = n9498_dest_is_safe_v[7];
  assign n9667_o = n9498_dest_is_safe_v[15:11];
  assign n9668_o = {n9667_o, n9593_o, n9588_o, n9583_o, n9666_o, n9578_o, n9573_o, n9568_o, n9665_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1582:163  */
  assign n9669_o = n9668_o[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1582:123  */
  assign n9670_o = n9664_o & n9669_o;
  assign n9671_o = n9498_source_is_safe_v[3];
  assign n9672_o = n9498_source_is_safe_v[7];
  assign n9673_o = n9498_source_is_safe_v[15:11];
  assign n9674_o = {n9673_o, n9548_o, n9543_o, n9538_o, n9672_o, n9533_o, n9528_o, n9523_o, n9671_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1583:96  */
  assign n9675_o = n9674_o[9];
  assign n9676_o = n9498_dest_is_safe_v[3];
  assign n9677_o = n9498_dest_is_safe_v[7];
  assign n9678_o = n9498_dest_is_safe_v[15:11];
  assign n9679_o = {n9678_o, n9593_o, n9588_o, n9583_o, n9677_o, n9578_o, n9573_o, n9568_o, n9676_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1583:151  */
  assign n9680_o = n9679_o[6];
  /* ../../HW/src/dp/dp_fetch.vhd:1583:115  */
  assign n9681_o = n9675_o & n9680_o;
  assign n9682_o = n9498_source_is_safe_v[3];
  assign n9683_o = n9498_source_is_safe_v[7];
  assign n9684_o = n9498_source_is_safe_v[15:11];
  assign n9685_o = {n9684_o, n9548_o, n9543_o, n9538_o, n9683_o, n9533_o, n9528_o, n9523_o, n9682_o, n9518_o, n9513_o, n9508_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1584:95  */
  assign n9686_o = n9685_o[10];
  assign n9687_o = n9498_dest_is_safe_v[3];
  assign n9688_o = n9498_dest_is_safe_v[7];
  assign n9689_o = n9498_dest_is_safe_v[15:11];
  assign n9690_o = {n9689_o, n9593_o, n9588_o, n9583_o, n9688_o, n9578_o, n9573_o, n9568_o, n9687_o, n9563_o, n9558_o, n9553_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1584:148  */
  assign n9691_o = n9690_o[10];
  /* ../../HW/src/dp/dp_fetch.vhd:1584:113  */
  assign n9692_o = n9686_o & n9691_o;
  assign n9693_o = {n9626_o, n9615_o, n9604_o};
  assign n9694_o = {n9659_o, n9648_o, n9637_o};
  assign n9695_o = {n9692_o, n9681_o, n9670_o};
  assign n9702_o = {n9518_o, n9513_o, n9508_o};
  assign n9703_o = {n9533_o, n9528_o, n9523_o};
  assign n9704_o = {n9548_o, n9543_o, n9538_o};
  assign n9711_o = {n9563_o, n9558_o, n9553_o};
  assign n9712_o = {n9578_o, n9573_o, n9568_o};
  assign n9713_o = {n9593_o, n9588_o, n9583_o};
  assign n9723_o = new_cmd_is_safe_r[3];
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9724_o = n9502_o ? 1'b0 : n9723_o;
  assign n9728_o = new_cmd_is_safe_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9729_o = n9502_o ? 1'b0 : n9728_o;
  assign n9733_o = new_cmd_is_safe_r[15:11];
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9734_o = n9502_o ? 5'b00000 : n9733_o;
  assign n9748_o = n9499_o[10:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1534:1  */
  assign n9749_o = ~n9502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9750_o = n9498_source_is_safe_v[10:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9751_o = n9749_o ? n9704_o : n9750_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in)
    n9752_q <= n9751_o;
  initial
    n9752_q = n9748_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9753_o = n9499_o[6:4];
  /* ../../HW/src/dp/dp_fetch.vhd:1534:1  */
  assign n9754_o = ~n9502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9755_o = n9498_source_is_safe_v[6:4];
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9756_o = n9754_o ? n9703_o : n9755_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in)
    n9757_q <= n9756_o;
  initial
    n9757_q = n9753_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9758_o = n9499_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1534:1  */
  assign n9759_o = ~n9502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9760_o = n9498_source_is_safe_v[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9761_o = n9759_o ? n9702_o : n9760_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in)
    n9762_q <= n9761_o;
  initial
    n9762_q = n9758_o;
  assign n9766_o = {5'bZ, n9752_q, 1'bZ, n9757_q, 1'bZ, n9762_q};
  assign n9767_o = n9500_o[10:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1534:1  */
  assign n9768_o = ~n9502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9769_o = n9498_dest_is_safe_v[10:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9770_o = n9768_o ? n9713_o : n9769_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in)
    n9771_q <= n9770_o;
  initial
    n9771_q = n9767_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9772_o = n9500_o[6:4];
  /* ../../HW/src/dp/dp_fetch.vhd:1534:1  */
  assign n9773_o = ~n9502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9774_o = n9498_dest_is_safe_v[6:4];
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9775_o = n9773_o ? n9712_o : n9774_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in)
    n9776_q <= n9775_o;
  initial
    n9776_q = n9772_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n9777_o = n9500_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1534:1  */
  assign n9778_o = ~n9502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9779_o = n9498_dest_is_safe_v[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  assign n9780_o = n9778_o ? n9711_o : n9779_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in)
    n9781_q <= n9780_o;
  initial
    n9781_q = n9777_o;
  assign n9785_o = {5'bZ, n9771_q, 1'bZ, n9776_q, 1'bZ, n9781_q};
  /* ../../HW/src/dp/dp_fetch.vhd:1590:13  */
  assign n9787_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1590:17  */
  assign n9788_o = n9787_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1590:24  */
  assign n9790_o = n9788_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1591:13  */
  assign n9791_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1591:17  */
  assign n9792_o = n9791_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1591:24  */
  assign n9794_o = n9792_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1590:48  */
  assign n9795_o = n9794_o & n9790_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1592:13  */
  assign n9796_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1592:17  */
  assign n9797_o = n9796_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1592:27  */
  assign n9799_o = n9797_o == 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1591:48  */
  assign n9800_o = n9799_o & n9795_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1594:13  */
  assign n9801_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1594:17  */
  assign n9802_o = n9801_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1594:28  */
  assign n9803_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1594:32  */
  assign n9804_o = n9803_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1594:20  */
  assign n9805_o = n9802_o != n9804_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1596:26  */
  assign n9806_o = orecs[3];
  /* ../../HW/src/dp/dp_fetch.vhd:1596:57  */
  assign n9807_o = ~n9806_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1596:71  */
  assign n9808_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1596:75  */
  assign n9809_o = n9808_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1596:87  */
  assign n9811_o = n9809_o != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1596:119  */
  assign n9812_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1596:123  */
  assign n9813_o = n9812_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1596:137  */
  assign n9815_o = n9813_o != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1596:110  */
  assign n9816_o = n9815_o & n9811_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1596:62  */
  assign n9817_o = n9807_o | n9816_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1597:26  */
  assign n9818_o = orecs[4];
  /* ../../HW/src/dp/dp_fetch.vhd:1597:53  */
  assign n9819_o = ~n9818_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1597:67  */
  assign n9820_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1597:71  */
  assign n9821_o = n9820_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1597:83  */
  assign n9823_o = n9821_o != 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:1597:111  */
  assign n9824_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1597:115  */
  assign n9825_o = n9824_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1597:129  */
  assign n9827_o = n9825_o != 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:1597:102  */
  assign n9828_o = n9827_o & n9823_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1597:58  */
  assign n9829_o = n9819_o | n9828_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1596:162  */
  assign n9830_o = n9829_o & n9817_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1598:26  */
  assign n9831_o = orecs[6];
  /* ../../HW/src/dp/dp_fetch.vhd:1598:52  */
  assign n9832_o = ~n9831_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1598:66  */
  assign n9833_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1598:70  */
  assign n9834_o = n9833_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1598:82  */
  assign n9836_o = n9834_o != 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:1598:109  */
  assign n9837_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1598:113  */
  assign n9838_o = n9837_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1598:127  */
  assign n9840_o = n9838_o != 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:1598:100  */
  assign n9841_o = n9840_o & n9836_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1598:57  */
  assign n9842_o = n9832_o | n9841_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1597:150  */
  assign n9843_o = n9842_o & n9830_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1594:36  */
  assign n9844_o = n9805_o | n9843_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1592:85  */
  assign n9845_o = n9844_o & n9800_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1589:21  */
  assign n9846_o = n9845_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1606:13  */
  assign n9851_o = pauses[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1606:16  */
  assign n9852_o = ~n9851_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1608:20  */
  assign n9853_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1609:22  */
  assign n9854_o = valids[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1612:22  */
  assign n9856_o = pauses[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1613:16  */
  assign n9857_o = pauses[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1613:19  */
  assign n9858_o = ~n9857_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1613:24  */
  assign n9859_o = outoforderok & n9858_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1615:20  */
  assign n9860_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1616:22  */
  assign n9861_o = valids[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1619:22  */
  assign n9863_o = pauses[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1621:20  */
  assign n9864_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1622:22  */
  assign n9865_o = valids[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1625:22  */
  assign n9867_o = pauses[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1613:4  */
  assign n9868_o = n9859_o ? n9860_o : n9864_o;
  assign n9869_o = {1'b0, rdreq};
  assign n9870_o = {rdreq, 1'b0};
  /* ../../HW/src/dp/dp_fetch.vhd:1613:4  */
  assign n9871_o = n9859_o ? n9870_o : n9869_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1613:4  */
  assign n9872_o = n9859_o ? n9861_o : n9865_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1613:4  */
  assign n9873_o = n9859_o ? n9863_o : n9867_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1606:4  */
  assign n9874_o = n9852_o ? n9853_o : n9868_o;
  assign n9875_o = {1'b0, rdreq};
  /* ../../HW/src/dp/dp_fetch.vhd:1606:4  */
  assign n9876_o = n9852_o ? n9875_o : n9871_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1606:4  */
  assign n9877_o = n9852_o ? n9854_o : n9872_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1606:4  */
  assign n9878_o = n9852_o ? n9856_o : n9873_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1641:10  */
  assign n9883_o = valids[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:17  */
  assign n9885_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:21  */
  assign n9886_o = n9885_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:28  */
  assign n9888_o = n9886_o != 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:63  */
  assign n9889_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:67  */
  assign n9890_o = n9889_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:103  */
  assign n9891_o = condition_vm0_busy_r | condition_vm1_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:77  */
  assign n9892_o = n9890_o & n9891_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:129  */
  assign n9894_o = n9892_o != 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:53  */
  assign n9895_o = n9894_o & n9888_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:17  */
  assign n9897_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:21  */
  assign n9898_o = n9897_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:28  */
  assign n9900_o = n9898_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:62  */
  assign n9901_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:66  */
  assign n9902_o = n9901_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:68  */
  assign n9903_o = ~n9902_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:52  */
  assign n9904_o = n9903_o & n9900_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:84  */
  assign n9905_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:88  */
  assign n9906_o = n9905_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:98  */
  assign n9907_o = n9906_o & condition_vm0_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:124  */
  assign n9909_o = n9907_o != 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:74  */
  assign n9910_o = n9909_o & n9904_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:17  */
  assign n9912_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:21  */
  assign n9913_o = n9912_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:28  */
  assign n9915_o = n9913_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:62  */
  assign n9916_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:66  */
  assign n9917_o = n9916_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:52  */
  assign n9918_o = n9917_o & n9915_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:84  */
  assign n9919_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:88  */
  assign n9920_o = n9919_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:98  */
  assign n9921_o = n9920_o & condition_vm1_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:124  */
  assign n9923_o = n9921_o != 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:74  */
  assign n9924_o = n9923_o & n9918_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:20  */
  assign n9926_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:24  */
  assign n9927_o = n9926_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:30  */
  assign n9929_o = n9927_o == 3'b100;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:60  */
  assign n9930_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:64  */
  assign n9931_o = n9930_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:66  */
  assign n9932_o = ~n9931_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:51  */
  assign n9933_o = n9932_o & n9929_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1654:9  */
  assign n9936_o = task_r ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1659:16  */
  assign n9937_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:20  */
  assign n9938_o = n9937_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:26  */
  assign n9940_o = n9938_o == 3'b100;
  /* ../../HW/src/dp/dp_fetch.vhd:1659:56  */
  assign n9941_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:60  */
  assign n9942_o = n9941_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:47  */
  assign n9943_o = n9942_o & n9940_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1662:9  */
  assign n9946_o = task_r ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1667:16  */
  assign n9947_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1667:20  */
  assign n9948_o = n9947_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1667:27  */
  assign n9950_o = n9948_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:22  */
  assign n9951_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:26  */
  assign n9952_o = n9951_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:39  */
  assign n9954_o = n9952_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:102  */
  assign n9955_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:106  */
  assign n9956_o = n9955_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:108  */
  assign n9957_o = n9956_o == task_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:93  */
  assign n9958_o = n9957_o & n9954_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1671:22  */
  assign n9959_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:26  */
  assign n9960_o = n9959_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:37  */
  assign n9962_o = n9960_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1671:100  */
  assign n9963_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:104  */
  assign n9964_o = n9963_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:106  */
  assign n9965_o = n9964_o == task_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1671:91  */
  assign n9966_o = n9965_o & n9962_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:120  */
  assign n9967_o = n9958_o | n9966_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1668:24  */
  assign n9968_o = n9967_o & task_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1678:64  */
  assign n9970_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:68  */
  assign n9971_o = n9970_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:100  */
  assign n9974_o = orecs[1619:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:104  */
  assign n9975_o = n9974_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:26  */
  assign n9980_o = ~n11043_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1668:10  */
  assign n9981_o = n9968_o ? 1'b1 : n9980_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1667:5  */
  assign n9983_o = n9950_o ? n9981_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1659:5  */
  assign n9984_o = n9943_o ? n9946_o : n9983_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:9  */
  assign n9985_o = n9933_o ? n9936_o : n9984_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:5  */
  assign n9986_o = n9924_o ? 1'b1 : n9985_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:5  */
  assign n9987_o = n9910_o ? 1'b1 : n9986_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:5  */
  assign n9988_o = n9895_o ? 1'b1 : n9987_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1642:5  */
  assign n9989_o = indication_full_r ? 1'b1 : n9988_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1641:1  */
  assign n9991_o = n9883_o ? n9989_o : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1641:10  */
  assign n9992_o = valids[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:17  */
  assign n9994_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:21  */
  assign n9995_o = n9994_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:28  */
  assign n9997_o = n9995_o != 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:63  */
  assign n9998_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:67  */
  assign n9999_o = n9998_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1644:103  */
  assign n10000_o = condition_vm0_busy_r | condition_vm1_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:77  */
  assign n10001_o = n9999_o & n10000_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:129  */
  assign n10003_o = n10001_o != 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:53  */
  assign n10004_o = n10003_o & n9997_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:17  */
  assign n10006_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:21  */
  assign n10007_o = n10006_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:28  */
  assign n10009_o = n10007_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:62  */
  assign n10010_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:66  */
  assign n10011_o = n10010_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:68  */
  assign n10012_o = ~n10011_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:52  */
  assign n10013_o = n10012_o & n10009_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:84  */
  assign n10014_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:88  */
  assign n10015_o = n10014_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1647:98  */
  assign n10016_o = n10015_o & condition_vm0_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:124  */
  assign n10018_o = n10016_o != 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:74  */
  assign n10019_o = n10018_o & n10013_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:17  */
  assign n10021_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:21  */
  assign n10022_o = n10021_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:28  */
  assign n10024_o = n10022_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:62  */
  assign n10025_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:66  */
  assign n10026_o = n10025_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:52  */
  assign n10027_o = n10026_o & n10024_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:84  */
  assign n10028_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:88  */
  assign n10029_o = n10028_o[6:3];
  /* ../../HW/src/dp/dp_fetch.vhd:1649:98  */
  assign n10030_o = n10029_o & condition_vm1_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:124  */
  assign n10032_o = n10030_o != 4'b0000;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:74  */
  assign n10033_o = n10032_o & n10027_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:20  */
  assign n10035_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:24  */
  assign n10036_o = n10035_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:30  */
  assign n10038_o = n10036_o == 3'b100;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:60  */
  assign n10039_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:64  */
  assign n10040_o = n10039_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1651:66  */
  assign n10041_o = ~n10040_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:51  */
  assign n10042_o = n10041_o & n10038_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1654:9  */
  assign n10045_o = task_r ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1659:16  */
  assign n10046_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:20  */
  assign n10047_o = n10046_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:26  */
  assign n10049_o = n10047_o == 3'b100;
  /* ../../HW/src/dp/dp_fetch.vhd:1659:56  */
  assign n10050_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:60  */
  assign n10051_o = n10050_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1659:47  */
  assign n10052_o = n10051_o & n10049_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1662:9  */
  assign n10055_o = task_r ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1667:16  */
  assign n10056_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1667:20  */
  assign n10057_o = n10056_o[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1667:27  */
  assign n10059_o = n10057_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:22  */
  assign n10060_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:26  */
  assign n10061_o = n10060_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:39  */
  assign n10063_o = n10061_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:102  */
  assign n10064_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:106  */
  assign n10065_o = n10064_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1670:108  */
  assign n10066_o = n10065_o == task_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:93  */
  assign n10067_o = n10066_o & n10063_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1671:22  */
  assign n10068_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:26  */
  assign n10069_o = n10068_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:37  */
  assign n10071_o = n10069_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1671:100  */
  assign n10072_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:104  */
  assign n10073_o = n10072_o[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1671:106  */
  assign n10074_o = n10073_o == task_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1671:91  */
  assign n10075_o = n10074_o & n10071_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1670:120  */
  assign n10076_o = n10067_o | n10075_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1668:24  */
  assign n10077_o = n10076_o & task_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1678:64  */
  assign n10079_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:68  */
  assign n10080_o = n10079_o[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:100  */
  assign n10083_o = orecs[3239:1620];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:104  */
  assign n10084_o = n10083_o[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:26  */
  assign n10089_o = ~n11070_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1668:10  */
  assign n10090_o = n10077_o ? 1'b1 : n10089_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1667:5  */
  assign n10092_o = n10059_o ? n10090_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1659:5  */
  assign n10093_o = n10052_o ? n10055_o : n10092_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1651:9  */
  assign n10094_o = n10042_o ? n10045_o : n10093_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1649:5  */
  assign n10095_o = n10033_o ? 1'b1 : n10094_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1647:5  */
  assign n10096_o = n10019_o ? 1'b1 : n10095_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1644:5  */
  assign n10097_o = n10004_o ? 1'b1 : n10096_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1642:5  */
  assign n10098_o = indication_full_r ? 1'b1 : n10097_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1641:1  */
  assign n10100_o = n9992_o ? n10098_o : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1696:10  */
  assign n10104_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1696:16  */
  assign n10106_o = n10104_o == 3'b110;
  /* ../../HW/src/dp/dp_fetch.vhd:1695:14  */
  assign n10107_o = n10106_o & ready;
  /* ../../HW/src/dp/dp_fetch.vhd:1697:10  */
  assign n10108_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1696:72  */
  assign n10109_o = n10108_o & n10107_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1695:1  */
  assign n10112_o = n10109_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1706:13  */
  assign n10116_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1713:47  */
  assign n10118_o = orec_generic[96:33];
  /* ../../HW/src/dp/dp_fetch.vhd:1716:29  */
  assign n10119_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1716:35  */
  assign n10121_o = n10119_o == 3'b111;
  /* ../../HW/src/dp/dp_fetch.vhd:1716:20  */
  assign n10122_o = n10121_o & ready;
  /* ../../HW/src/dp/dp_fetch.vhd:1716:95  */
  assign n10123_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1716:86  */
  assign n10124_o = n10123_o & n10122_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1716:7  */
  assign n10127_o = n10124_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1733:11  */
  assign n10144_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1733:17  */
  assign n10146_o = n10144_o == 3'b100;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:14  */
  assign n10147_o = n10146_o & ready;
  /* ../../HW/src/dp/dp_fetch.vhd:1733:81  */
  assign n10148_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1733:83  */
  assign n10149_o = ~n10148_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1733:71  */
  assign n10150_o = n10149_o & n10147_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1734:10  */
  assign n10151_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1733:89  */
  assign n10152_o = n10151_o & n10150_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1738:42  */
  assign n10153_o = orec_generic[18:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1740:46  */
  assign n10154_o = orec_generic[23:19];
  /* ../../HW/src/dp/dp_fetch.vhd:1742:40  */
  assign n10155_o = orec_generic[24];
  /* ../../HW/src/dp/dp_fetch.vhd:1744:140  */
  assign n10156_o = orec_generic[26:25];
  /* ../../HW/src/dp/dp_fetch.vhd:1746:40  */
  assign n10157_o = orec_generic[30:27];
  /* ../../HW/src/dp/dp_fetch.vhd:1748:42  */
  assign n10158_o = orec_generic[32:31];
  /* ../../HW/src/dp/dp_fetch.vhd:1751:118  */
  assign n10159_o = orec_generic[45:33];
  /* ../../HW/src/dp/dp_fetch.vhd:1751:118  */
  assign n10160_o = orec_generic[77:65];
  /* ../../HW/src/dp/dp_fetch.vhd:1754:11  */
  assign n10161_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1754:17  */
  assign n10163_o = n10161_o == 3'b100;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:17  */
  assign n10164_o = n10163_o & ready;
  /* ../../HW/src/dp/dp_fetch.vhd:1754:81  */
  assign n10165_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1754:71  */
  assign n10166_o = n10165_o & n10164_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1755:10  */
  assign n10167_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1754:89  */
  assign n10168_o = n10167_o & n10166_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1759:42  */
  assign n10169_o = orec_generic[18:8];
  /* ../../HW/src/dp/dp_fetch.vhd:1761:46  */
  assign n10170_o = orec_generic[23:19];
  /* ../../HW/src/dp/dp_fetch.vhd:1763:40  */
  assign n10171_o = orec_generic[24];
  /* ../../HW/src/dp/dp_fetch.vhd:1765:140  */
  assign n10172_o = orec_generic[26:25];
  /* ../../HW/src/dp/dp_fetch.vhd:1767:40  */
  assign n10173_o = orec_generic[30:27];
  /* ../../HW/src/dp/dp_fetch.vhd:1769:42  */
  assign n10174_o = orec_generic[32:31];
  /* ../../HW/src/dp/dp_fetch.vhd:1772:117  */
  assign n10175_o = orec_generic[45:33];
  /* ../../HW/src/dp/dp_fetch.vhd:1772:117  */
  assign n10176_o = orec_generic[77:65];
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10178_o = n10168_o ? n10169_o : 11'b00000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10180_o = n10168_o ? n10170_o : 5'b11111;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10182_o = n10168_o ? n10173_o : 4'b1111;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10184_o = n10168_o ? n10174_o : 2'b00;
  assign n10185_o = {n10172_o, n10176_o, n10175_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10187_o = n10168_o ? n10185_o : 28'b0000000000000000000000000000;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10189_o = n10168_o ? n10171_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10192_o = n10168_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1753:1  */
  assign n10195_o = n10168_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10198_o = n10152_o ? n10153_o : n10178_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10199_o = n10152_o ? n10154_o : n10180_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10200_o = n10152_o ? n10157_o : n10182_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10201_o = n10152_o ? n10158_o : n10184_o;
  assign n10202_o = {n10156_o, n10160_o, n10159_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10203_o = n10152_o ? n10202_o : n10187_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10204_o = n10152_o ? n10155_o : n10189_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10206_o = n10152_o ? 1'b1 : n10192_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1732:1  */
  assign n10208_o = n10152_o ? 1'b0 : n10195_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1795:12  */
  assign n10214_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1795:19  */
  assign n10216_o = n10214_o == 3'b001;
  /* ../../HW/src/dp/dp_fetch.vhd:1796:16  */
  assign n10217_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1795:4  */
  assign n10219_o = n10216_o ? n10217_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1794:1  */
  assign n10221_o = ready ? n10219_o : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1807:17  */
  assign n10225_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1811:34  */
  assign n10227_o = ~pause;
  /* ../../HW/src/dp/dp_fetch.vhd:1811:25  */
  assign n10228_o = n10227_o & ready;
  /* ../../HW/src/dp/dp_fetch.vhd:1812:23  */
  assign n10229_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1812:30  */
  assign n10231_o = n10229_o == 3'b010;
  /* ../../HW/src/dp/dp_fetch.vhd:1814:26  */
  assign n10232_o = orec[2:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1814:33  */
  assign n10234_o = n10232_o == 3'b011;
  /* ../../HW/src/dp/dp_fetch.vhd:1814:15  */
  assign n10236_o = n10234_o ? 1'b0 : log_enable_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1812:15  */
  assign n10238_o = n10231_o ? 1'b1 : n10236_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1824:17  */
  assign n10246_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1836:22  */
  assign n10248_o = ~task_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1846:13  */
  assign n10250_o = task2 ? 1'b0 : task_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1836:13  */
  assign n10258_o = n10248_o ? \task  : n10250_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1862:17  */
  assign n10292_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1870:20  */
  assign n10294_o = ~wreq2;
  /* ../../HW/src/dp/dp_fetch.vhd:1873:29  */
  assign n10295_o = ~ready_which;
  /* ../../HW/src/dp/dp_fetch.vhd:1876:52  */
  assign n10297_o = instruction[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1877:48  */
  assign n10298_o = instruction[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1878:50  */
  assign n10299_o = instruction[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1882:52  */
  assign n10301_o = instruction[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:1883:48  */
  assign n10302_o = instruction[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1884:50  */
  assign n10303_o = instruction[1565:1564];
  assign n10304_o = {wreq2, 1'b0};
  assign n10305_o = {1'b0, wreq2};
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10306_o = n10295_o ? n10305_o : n10304_o;
  assign n10307_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10308_o = n10295_o ? n10297_o : n10307_o;
  assign n10309_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10310_o = n10295_o ? n10309_o : n10301_o;
  assign n10311_o = source_vm_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10312_o = n10295_o ? n10298_o : n10311_o;
  assign n10313_o = source_vm_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10314_o = n10295_o ? n10313_o : n10302_o;
  assign n10315_o = dest_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10316_o = n10295_o ? n10299_o : n10315_o;
  assign n10317_o = dest_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1873:15  */
  assign n10318_o = n10295_o ? n10317_o : n10303_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1870:12  */
  assign n10320_o = n10294_o ? 2'b00 : n10306_o;
  assign n10321_o = {n10310_o, n10308_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1870:12  */
  assign n10322_o = n10294_o ? source_bus_id_r : n10321_o;
  assign n10323_o = {n10314_o, n10312_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1870:12  */
  assign n10324_o = n10294_o ? source_vm_r : n10323_o;
  assign n10325_o = {n10318_o, n10316_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1870:12  */
  assign n10326_o = n10294_o ? dest_bus_id_r : n10325_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1908:16  */
  assign n10356_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1928:42  */
  assign n10359_o = $unsigned(indication_wrusedw) >= $unsigned(8'b11110111);
  /* ../../HW/src/dp/dp_fetch.vhd:1928:10  */
  assign n10362_o = n10359_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1934:33  */
  assign n10363_o = pcore_sink_counter_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1934:58  */
  assign n10364_o = pcore_sink_counter_in[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1934:36  */
  assign n10365_o = n10363_o == n10364_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1934:10  */
  assign n10368_o = n10365_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1939:33  */
  assign n10369_o = pcore_sink_counter_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1939:58  */
  assign n10370_o = pcore_sink_counter_in[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1939:36  */
  assign n10371_o = n10369_o == n10370_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1939:10  */
  assign n10374_o = n10371_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1944:32  */
  assign n10375_o = sram_sink_counter_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1944:56  */
  assign n10376_o = sram_sink_counter_in[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1944:35  */
  assign n10377_o = n10375_o == n10376_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1944:10  */
  assign n10380_o = n10377_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1949:32  */
  assign n10381_o = sram_sink_counter_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1949:56  */
  assign n10382_o = sram_sink_counter_in[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1949:35  */
  assign n10383_o = n10381_o == n10382_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1949:10  */
  assign n10386_o = n10383_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1954:31  */
  assign n10387_o = ddr_sink_counter_r == ddr_sink_counter_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1954:10  */
  assign n10390_o = n10387_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1961:33  */
  assign n10392_o = instruction_valid_r != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1962:38  */
  assign n10393_o = instruction_r[1597:1574];
  /* ../../HW/src/dp/dp_fetch.vhd:1963:30  */
  assign n10394_o = instruction_r[1563:788];
  /* ../../HW/src/dp/dp_fetch.vhd:1963:35  */
  assign n10395_o = n10394_o[673];
  /* ../../HW/src/dp/dp_fetch.vhd:1963:74  */
  assign n10396_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1963:86  */
  assign n10398_o = n10396_o != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1963:56  */
  assign n10399_o = n10398_o & n10395_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1964:35  */
  assign n10401_o = n10393_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_fetch.vhd:1963:13  */
  assign n10402_o = n10399_o ? n10401_o : n10393_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1966:30  */
  assign n10403_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1966:41  */
  assign n10405_o = n10403_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1967:33  */
  assign n10406_o = instruction_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1967:35  */
  assign n10407_o = ~n10406_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1968:66  */
  assign n10408_o = pcore_sink_counter_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1968:69  */
  assign n10409_o = n10408_o + n10402_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1971:66  */
  assign n10411_o = pcore_sink_counter_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1971:69  */
  assign n10412_o = n10411_o + n10402_o;
  assign n10414_o = pcore_sink_counter_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1967:16  */
  assign n10415_o = n10407_o ? n10409_o : n10414_o;
  assign n10416_o = pcore_sink_counter_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1967:16  */
  assign n10417_o = n10407_o ? n10416_o : n10412_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1967:16  */
  assign n10418_o = n10407_o ? 1'b1 : n10368_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1967:16  */
  assign n10419_o = n10407_o ? n10374_o : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1974:36  */
  assign n10420_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1974:47  */
  assign n10422_o = n10420_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:1975:36  */
  assign n10423_o = instruction_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1975:38  */
  assign n10424_o = ~n10423_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1976:67  */
  assign n10425_o = sram_sink_counter_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1976:70  */
  assign n10426_o = n10425_o + n10402_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1979:67  */
  assign n10428_o = sram_sink_counter_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1979:70  */
  assign n10429_o = n10428_o + n10402_o;
  assign n10431_o = sram_sink_counter_r[23:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1975:19  */
  assign n10432_o = n10424_o ? n10426_o : n10431_o;
  assign n10433_o = sram_sink_counter_r[47:24];
  /* ../../HW/src/dp/dp_fetch.vhd:1975:19  */
  assign n10434_o = n10424_o ? n10433_o : n10429_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1975:19  */
  assign n10435_o = n10424_o ? 1'b1 : n10380_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1975:19  */
  assign n10436_o = n10424_o ? n10386_o : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1983:59  */
  assign n10437_o = ddr_sink_counter_r + n10402_o;
  assign n10438_o = {n10434_o, n10432_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1974:16  */
  assign n10439_o = n10422_o ? n10438_o : sram_sink_counter_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1974:16  */
  assign n10440_o = n10422_o ? ddr_sink_counter_r : n10437_o;
  assign n10441_o = {n10436_o, n10435_o};
  assign n10442_o = {n10386_o, n10380_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1974:16  */
  assign n10443_o = n10422_o ? n10441_o : n10442_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1974:16  */
  assign n10445_o = n10422_o ? n10390_o : 1'b1;
  assign n10446_o = {n10417_o, n10415_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1966:13  */
  assign n10448_o = n10405_o ? sram_sink_counter_r : n10439_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1966:13  */
  assign n10449_o = n10405_o ? ddr_sink_counter_r : n10440_o;
  assign n10450_o = {n10419_o, n10418_o};
  assign n10451_o = {n10374_o, n10368_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1966:13  */
  assign n10452_o = n10405_o ? n10450_o : n10451_o;
  assign n10453_o = {n10386_o, n10380_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1966:13  */
  assign n10454_o = n10405_o ? n10453_o : n10443_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1966:13  */
  assign n10455_o = n10405_o ? n10390_o : n10445_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1961:10  */
  assign n10456_o = n10405_o & n10392_o;
  assign n10459_o = {n10374_o, n10368_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1961:10  */
  assign n10460_o = n10392_o ? n10452_o : n10459_o;
  assign n10461_o = {n10386_o, n10380_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1961:10  */
  assign n10462_o = n10392_o ? n10454_o : n10461_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1961:10  */
  assign n10463_o = n10392_o ? n10455_o : n10390_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1989:22  */
  assign n10466_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:1990:21  */
  assign n10467_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1990:32  */
  assign n10469_o = n10467_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1989:29  */
  assign n10470_o = n10469_o & n10466_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1990:95  */
  assign n10471_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1990:97  */
  assign n10472_o = ~n10471_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1990:86  */
  assign n10473_o = n10472_o & n10470_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1992:39  */
  assign n10476_o = instruction_valid_r != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1993:33  */
  assign n10477_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:1993:44  */
  assign n10479_o = n10477_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:1992:47  */
  assign n10480_o = n10479_o & n10476_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1994:33  */
  assign n10481_o = instruction_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1994:35  */
  assign n10482_o = ~n10481_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1993:98  */
  assign n10483_o = n10482_o & n10480_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1996:36  */
  assign n10485_o = pcore_sink_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1996:39  */
  assign n10486_o = ~n10485_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1996:13  */
  assign n10489_o = n10486_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:1992:13  */
  assign n10490_o = n10483_o ? 1'b1 : n10489_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1989:13  */
  assign n10491_o = n10473_o ? 1'b1 : n10490_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2004:22  */
  assign n10493_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2004:38  */
  assign n10494_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2004:49  */
  assign n10496_o = n10494_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2004:29  */
  assign n10497_o = n10496_o & n10493_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2004:112  */
  assign n10498_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2004:103  */
  assign n10499_o = n10498_o & n10497_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2006:39  */
  assign n10502_o = instruction_valid_r != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2007:30  */
  assign n10503_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2007:41  */
  assign n10505_o = n10503_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2006:47  */
  assign n10506_o = n10505_o & n10502_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2008:30  */
  assign n10507_o = instruction_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2007:95  */
  assign n10508_o = n10507_o & n10506_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2010:36  */
  assign n10510_o = pcore_sink_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2010:39  */
  assign n10511_o = ~n10510_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2010:13  */
  assign n10514_o = n10511_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:2006:13  */
  assign n10515_o = n10508_o ? 1'b1 : n10514_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2004:13  */
  assign n10516_o = n10499_o ? 1'b1 : n10515_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2018:22  */
  assign n10518_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2018:38  */
  assign n10519_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2018:49  */
  assign n10521_o = n10519_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2018:29  */
  assign n10522_o = n10521_o & n10518_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2018:108  */
  assign n10523_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2018:110  */
  assign n10524_o = ~n10523_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2018:99  */
  assign n10525_o = n10524_o & n10522_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2020:39  */
  assign n10528_o = instruction_valid_r != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2020:65  */
  assign n10529_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2020:76  */
  assign n10531_o = n10529_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2020:47  */
  assign n10532_o = n10531_o & n10528_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2020:135  */
  assign n10533_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2020:137  */
  assign n10534_o = ~n10533_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2020:126  */
  assign n10535_o = n10534_o & n10532_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2022:35  */
  assign n10537_o = sram_sink_busy_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2022:38  */
  assign n10538_o = ~n10537_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2022:13  */
  assign n10541_o = n10538_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:2020:13  */
  assign n10542_o = n10535_o ? 1'b1 : n10541_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2018:13  */
  assign n10543_o = n10525_o ? 1'b1 : n10542_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2028:22  */
  assign n10545_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2028:38  */
  assign n10546_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2028:49  */
  assign n10548_o = n10546_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2028:29  */
  assign n10549_o = n10548_o & n10545_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2028:108  */
  assign n10550_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2028:99  */
  assign n10551_o = n10550_o & n10549_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2030:39  */
  assign n10554_o = instruction_valid_r != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2030:65  */
  assign n10555_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2030:76  */
  assign n10557_o = n10555_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2030:47  */
  assign n10558_o = n10557_o & n10554_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2030:135  */
  assign n10559_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2030:126  */
  assign n10560_o = n10559_o & n10558_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2032:35  */
  assign n10562_o = sram_sink_busy_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2032:38  */
  assign n10563_o = ~n10562_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2032:13  */
  assign n10566_o = n10563_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:2030:13  */
  assign n10567_o = n10560_o ? 1'b1 : n10566_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2028:13  */
  assign n10568_o = n10551_o ? 1'b1 : n10567_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2040:22  */
  assign n10570_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2040:38  */
  assign n10571_o = orec[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2040:49  */
  assign n10573_o = n10571_o == 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:2040:29  */
  assign n10574_o = n10573_o & n10570_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2042:39  */
  assign n10576_o = instruction_valid_r != 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2042:65  */
  assign n10577_o = instruction_r[1565:1564];
  /* ../../HW/src/dp/dp_fetch.vhd:2042:76  */
  assign n10579_o = n10577_o == 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:2042:47  */
  assign n10580_o = n10579_o & n10576_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2044:34  */
  assign n10581_o = ~ddr_sink_busy_r;
  /* ../../HW/src/dp/dp_fetch.vhd:2044:57  */
  assign n10582_o = ~ddr_tx_busy_in;
  /* ../../HW/src/dp/dp_fetch.vhd:2044:39  */
  assign n10583_o = n10582_o & n10581_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2044:13  */
  assign n10586_o = n10583_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_fetch.vhd:2042:13  */
  assign n10588_o = n10580_o ? 1'b1 : n10586_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2040:13  */
  assign n10590_o = n10574_o ? 1'b1 : n10588_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:32  */
  assign n10591_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:2056:35  */
  assign n10593_o = n10591_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:104  */
  assign n10594_o = source_vm_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2056:107  */
  assign n10595_o = ~n10594_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:89  */
  assign n10596_o = n10595_o & n10593_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:122  */
  assign n10597_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2056:125  */
  assign n10598_o = ~n10597_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:112  */
  assign n10599_o = n10598_o & n10596_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2057:32  */
  assign n10600_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:2057:35  */
  assign n10602_o = n10600_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2057:104  */
  assign n10603_o = source_vm_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2057:107  */
  assign n10604_o = ~n10603_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2057:89  */
  assign n10605_o = n10604_o & n10602_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2057:122  */
  assign n10606_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2057:125  */
  assign n10607_o = ~n10606_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2057:112  */
  assign n10608_o = n10607_o & n10605_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:132  */
  assign n10609_o = n10599_o | n10608_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2058:41  */
  assign n10610_o = pcore_read_pending_p0_in[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2057:132  */
  assign n10611_o = n10609_o | n10610_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2059:40  */
  assign n10612_o = sram_read_pending_p0_in[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2058:69  */
  assign n10613_o = n10611_o | n10612_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2060:33  */
  assign n10614_o = ddr_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2059:68  */
  assign n10615_o = n10613_o | n10614_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2056:13  */
  assign n10618_o = n10615_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2066:32  */
  assign n10619_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:2066:35  */
  assign n10621_o = n10619_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2066:104  */
  assign n10622_o = source_vm_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2066:89  */
  assign n10623_o = n10622_o & n10621_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2066:122  */
  assign n10624_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2066:125  */
  assign n10625_o = ~n10624_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2066:112  */
  assign n10626_o = n10625_o & n10623_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2067:32  */
  assign n10627_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:2067:35  */
  assign n10629_o = n10627_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2067:104  */
  assign n10630_o = source_vm_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2067:89  */
  assign n10631_o = n10630_o & n10629_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2067:122  */
  assign n10632_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2067:125  */
  assign n10633_o = ~n10632_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2067:112  */
  assign n10634_o = n10633_o & n10631_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2066:132  */
  assign n10635_o = n10626_o | n10634_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2068:41  */
  assign n10636_o = pcore_read_pending_p1_in[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2067:132  */
  assign n10637_o = n10635_o | n10636_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2069:40  */
  assign n10638_o = sram_read_pending_p1_in[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2068:69  */
  assign n10639_o = n10637_o | n10638_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2070:33  */
  assign n10640_o = ddr_read_pending[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2069:68  */
  assign n10641_o = n10639_o | n10640_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2066:13  */
  assign n10644_o = n10641_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:32  */
  assign n10645_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:2078:35  */
  assign n10647_o = n10645_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:100  */
  assign n10648_o = source_vm_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2078:103  */
  assign n10649_o = ~n10648_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:85  */
  assign n10650_o = n10649_o & n10647_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:118  */
  assign n10651_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2078:121  */
  assign n10652_o = ~n10651_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:108  */
  assign n10653_o = n10652_o & n10650_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2079:32  */
  assign n10654_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:2079:35  */
  assign n10656_o = n10654_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2079:100  */
  assign n10657_o = source_vm_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2079:103  */
  assign n10658_o = ~n10657_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2079:85  */
  assign n10659_o = n10658_o & n10656_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2079:118  */
  assign n10660_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2079:121  */
  assign n10661_o = ~n10660_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2079:108  */
  assign n10662_o = n10661_o & n10659_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:128  */
  assign n10663_o = n10653_o | n10662_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2080:41  */
  assign n10664_o = pcore_read_pending_p0_in[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2079:128  */
  assign n10665_o = n10663_o | n10664_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2081:40  */
  assign n10666_o = sram_read_pending_p0_in[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2080:65  */
  assign n10667_o = n10665_o | n10666_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2082:33  */
  assign n10668_o = ddr_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2081:64  */
  assign n10669_o = n10667_o | n10668_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2078:13  */
  assign n10672_o = n10669_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2088:32  */
  assign n10673_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:2088:35  */
  assign n10675_o = n10673_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2088:100  */
  assign n10676_o = source_vm_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2088:85  */
  assign n10677_o = n10676_o & n10675_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2088:118  */
  assign n10678_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2088:121  */
  assign n10679_o = ~n10678_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2088:108  */
  assign n10680_o = n10679_o & n10677_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2089:32  */
  assign n10681_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:2089:35  */
  assign n10683_o = n10681_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2089:100  */
  assign n10684_o = source_vm_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2089:85  */
  assign n10685_o = n10684_o & n10683_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2089:118  */
  assign n10686_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2089:121  */
  assign n10687_o = ~n10686_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2089:108  */
  assign n10688_o = n10687_o & n10685_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2088:128  */
  assign n10689_o = n10680_o | n10688_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2090:41  */
  assign n10690_o = pcore_read_pending_p1_in[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2089:128  */
  assign n10691_o = n10689_o | n10690_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2091:40  */
  assign n10692_o = sram_read_pending_p1_in[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2090:65  */
  assign n10693_o = n10691_o | n10692_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2092:33  */
  assign n10694_o = ddr_read_pending[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2091:64  */
  assign n10695_o = n10693_o | n10694_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2088:13  */
  assign n10698_o = n10695_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2100:32  */
  assign n10699_o = source_bus_id_r[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:2100:35  */
  assign n10701_o = n10699_o == 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:2100:94  */
  assign n10702_o = avail[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2100:97  */
  assign n10703_o = ~n10702_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2100:84  */
  assign n10704_o = n10703_o & n10701_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2101:32  */
  assign n10705_o = source_bus_id_r[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:2101:35  */
  assign n10707_o = n10705_o == 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:2101:94  */
  assign n10708_o = avail[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2101:97  */
  assign n10709_o = ~n10708_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2101:84  */
  assign n10710_o = n10709_o & n10707_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2100:104  */
  assign n10711_o = n10704_o | n10710_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2102:35  */
  assign n10712_o = pcore_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:2101:104  */
  assign n10713_o = n10711_o | n10712_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2103:34  */
  assign n10714_o = sram_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:2102:58  */
  assign n10715_o = n10713_o | n10714_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2104:33  */
  assign n10716_o = ddr_read_pending[2];
  /* ../../HW/src/dp/dp_fetch.vhd:2103:57  */
  assign n10717_o = n10715_o | n10716_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2100:13  */
  assign n10720_o = n10717_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2112:22  */
  assign n10722_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2112:38  */
  assign n10723_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:2112:51  */
  assign n10725_o = n10723_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2112:29  */
  assign n10726_o = n10725_o & n10722_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2113:21  */
  assign n10727_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2113:23  */
  assign n10728_o = ~n10727_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2112:105  */
  assign n10729_o = n10728_o & n10726_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2112:13  */
  assign n10731_o = n10729_o ? 1'b1 : n10618_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2116:22  */
  assign n10733_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2116:38  */
  assign n10734_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:2116:51  */
  assign n10736_o = n10734_o == 2'b00;
  /* ../../HW/src/dp/dp_fetch.vhd:2116:29  */
  assign n10737_o = n10736_o & n10733_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2117:21  */
  assign n10738_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2116:105  */
  assign n10739_o = n10738_o & n10737_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2116:13  */
  assign n10741_o = n10739_o ? 1'b1 : n10644_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2121:22  */
  assign n10743_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2121:38  */
  assign n10744_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:2121:51  */
  assign n10746_o = n10744_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2121:29  */
  assign n10747_o = n10746_o & n10743_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2121:110  */
  assign n10748_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2121:112  */
  assign n10749_o = ~n10748_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2121:101  */
  assign n10750_o = n10749_o & n10747_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2121:13  */
  assign n10752_o = n10750_o ? 1'b1 : n10672_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2125:22  */
  assign n10754_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2125:38  */
  assign n10755_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:2125:51  */
  assign n10757_o = n10755_o == 2'b01;
  /* ../../HW/src/dp/dp_fetch.vhd:2125:29  */
  assign n10758_o = n10757_o & n10754_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2125:110  */
  assign n10759_o = orec[7];
  /* ../../HW/src/dp/dp_fetch.vhd:2125:101  */
  assign n10760_o = n10759_o & n10758_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2125:13  */
  assign n10762_o = n10760_o ? 1'b1 : n10698_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2129:22  */
  assign n10764_o = wreq2 != 1'b0;
  /* ../../HW/src/dp/dp_fetch.vhd:2129:38  */
  assign n10765_o = orec[785:784];
  /* ../../HW/src/dp/dp_fetch.vhd:2129:51  */
  assign n10767_o = n10765_o == 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:2129:29  */
  assign n10768_o = n10767_o & n10764_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2129:13  */
  assign n10770_o = n10768_o ? 1'b1 : n10720_o;
  assign n10771_o = {n10741_o, n10731_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2135:87  */
  assign n10772_o = n10771_o[0];
  assign n10773_o = {n10516_o, n10491_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2135:111  */
  assign n10774_o = n10773_o[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2135:91  */
  assign n10775_o = n10772_o | n10774_o;
  assign n10776_o = {n10762_o, n10752_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2136:82  */
  assign n10777_o = n10776_o[0];
  assign n10778_o = {n10568_o, n10543_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2136:105  */
  assign n10779_o = n10778_o[0];
  /* ../../HW/src/dp/dp_fetch.vhd:2136:86  */
  assign n10780_o = n10777_o | n10779_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2137:81  */
  assign n10781_o = n10770_o | n10590_o;
  assign n10782_o = {n10741_o, n10731_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2139:87  */
  assign n10783_o = n10782_o[1];
  assign n10784_o = {n10516_o, n10491_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2139:111  */
  assign n10785_o = n10784_o[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2139:91  */
  assign n10786_o = n10783_o | n10785_o;
  assign n10787_o = {n10762_o, n10752_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2140:82  */
  assign n10788_o = n10787_o[1];
  assign n10789_o = {n10568_o, n10543_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2140:105  */
  assign n10790_o = n10789_o[1];
  /* ../../HW/src/dp/dp_fetch.vhd:2140:86  */
  assign n10791_o = n10788_o | n10790_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2141:81  */
  assign n10792_o = n10770_o | n10590_o;
  assign n10793_o = {n10516_o, n10491_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2143:54  */
  assign n10794_o = n10793_o[0];
  assign n10795_o = {n10516_o, n10491_o};
  /* ../../HW/src/dp/dp_fetch.vhd:2144:54  */
  assign n10796_o = n10795_o[1];
  assign n10797_o = {n10568_o, n10543_o};
  assign n10798_o = {n10741_o, n10731_o};
  assign n10799_o = {n10762_o, n10752_o};
  assign n10803_o = {n10796_o, n10794_o};
  assign n10811_o = {n10780_o, n10775_o};
  assign n10816_o = {n10791_o, n10786_o};
  assign n10858_o = condition_vm0_busy_r[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n10859_o = n10356_o ? 1'b0 : n10858_o;
  assign n10865_o = condition_vm1_busy_r[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n10866_o = n10356_o ? 1'b0 : n10865_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2159:16  */
  assign n10908_o = ~reset_in;
  /* ../../HW/src/dp/dp_fetch.vhd:2164:34  */
  assign n10911_o = log_time_r + 32'b00000000000000000000000000000001;
  /* ../../HW/src/dp/dp_fetch.vhd:2165:40  */
  assign n10912_o = log_write[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:2165:71  */
  assign n10914_o = n10912_o != 2'b10;
  /* ../../HW/src/dp/dp_fetch.vhd:2165:27  */
  assign n10915_o = n10914_o & log_wrreq;
  assign n10924_o = {n8761_o, n8589_o};
  assign n10925_o = {n8859_o, n8850_o};
  assign n10926_o = {fifo_i_n7934, fifo_i_n7933};
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  assign n10927_o = n10456_o ? n10446_o : pcore_sink_counter_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10928_q <= 48'b000000000000000000000000000000000000000000000000;
    else
      n10928_q <= n10927_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  assign n10929_o = n10392_o ? n10448_o : sram_sink_counter_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10930_q <= 48'b000000000000000000000000000000000000000000000000;
    else
      n10930_q <= n10929_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  assign n10931_o = n10392_o ? n10449_o : ddr_sink_counter_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10932_q <= 24'b000000000000000000000000;
    else
      n10932_q <= n10931_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10933_q <= 2'b00;
    else
      n10933_q <= n10803_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10934_q <= 2'b00;
    else
      n10934_q <= n10797_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10935_q <= 1'b0;
    else
      n10935_q <= n10590_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10936_q <= 2'b00;
    else
      n10936_q <= n10798_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10937_q <= 2'b00;
    else
      n10937_q <= n10799_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10938_q <= 1'b0;
    else
      n10938_q <= n10770_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1810:9  */
  assign n10939_o = n10228_o ? n10238_o : log_enable_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1810:9  */
  always @(posedge clock_in or posedge n10225_o)
    if (n10225_o)
      n10940_q <= 1'b0;
    else
      n10940_q <= n10939_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1712:4  */
  always @(posedge clock_in or posedge n10116_o)
    if (n10116_o)
      n10941_q <= 1'b0;
    else
      n10941_q <= n10127_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1712:4  */
  always @(posedge clock_in or posedge n10116_o)
    if (n10116_o)
      n10942_q <= 1'b0;
    else
      n10942_q <= print_indication_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1712:4  */
  always @(posedge clock_in or posedge n10116_o)
    if (n10116_o)
      n10943_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n10943_q <= n10118_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1712:4  */
  always @(posedge clock_in or posedge n10116_o)
    if (n10116_o)
      n10944_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n10944_q <= print_param_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10945_q <= 1'b0;
    else
      n10945_q <= n10362_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  assign n10946_o = bus_write_r ? n9454_o : indication_parm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10947_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n10947_q <= n10946_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  assign n10948_o = n9009_o ? n8954_o : indication_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  always @(posedge clock_in or posedge n8947_o)
    if (n8947_o)
      n10949_q <= 32'b00000000000000000000000000000000;
    else
      n10949_q <= n10948_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  assign n10950_o = n9010_o ? 1'b0 : indication_sync_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  always @(posedge clock_in or posedge n8947_o)
    if (n8947_o)
      n10951_q <= 1'b0;
    else
      n10951_q <= n10950_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  assign n10952_o = n8951_o ? n9005_o : bus_readdata_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  always @(posedge clock_in or posedge n8947_o)
    if (n8947_o)
      n10953_q <= 32'b00000000000000000000000000000000;
    else
      n10953_q <= n10952_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in or posedge n10292_o)
    if (n10292_o)
      n10954_q <= 2'b00;
    else
      n10954_q <= n10320_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in or posedge n10292_o)
    if (n10292_o)
      n10955_q <= 2'b00;
    else
      n10955_q <= instruction_valid_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1860:1  */
  assign n10956_o = ~n10292_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  assign n10957_o = n10956_o ? instruction : instruction_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in)
    n10958_q <= n10957_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1860:1  */
  assign n10959_o = ~n10292_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  assign n10960_o = n10959_o ? instruction_r : instruction_rr;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in)
    n10961_q <= n10960_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2163:7  */
  assign n10962_o = n10915_o ? log_write : log_status_last_r;
  /* ../../HW/src/dp/dp_fetch.vhd:2163:7  */
  always @(posedge clock_in or posedge n10908_o)
    if (n10908_o)
      n10963_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n10963_q <= n10962_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  assign n10964_o = n8951_o ? n9006_o : log_readtime_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  always @(posedge clock_in or posedge n8947_o)
    if (n8947_o)
      n10965_q <= 32'b00000000000000000000000000000000;
    else
      n10965_q <= n10964_o;
  /* ../../HW/src/dp/dp_fetch.vhd:2163:7  */
  always @(posedge clock_in or posedge n10908_o)
    if (n10908_o)
      n10966_q <= 32'b00000000000000000000000000000000;
    else
      n10966_q <= n10911_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10968_q <= 1'b0;
    else
      n10968_q <= n9463_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  assign n10969_o = n9456_o ? n9318_o : load_busid_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10970_q <= 4'b0000;
    else
      n10970_q <= n10969_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in or posedge n10292_o)
    if (n10292_o)
      n10971_q <= 4'b0000;
    else
      n10971_q <= n10322_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in or posedge n10292_o)
    if (n10292_o)
      n10972_q <= 2'b00;
    else
      n10972_q <= n10324_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1869:9  */
  always @(posedge clock_in or posedge n10292_o)
    if (n10292_o)
      n10973_q <= 4'b0000;
    else
      n10973_q <= n10326_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in or posedge n9502_o)
    if (n9502_o)
      n10974_q <= 3'b000;
    else
      n10974_q <= n9695_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in or posedge n9502_o)
    if (n9502_o)
      n10975_q <= 3'b000;
    else
      n10975_q <= n9694_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1541:4  */
  always @(posedge clock_in or posedge n9502_o)
    if (n9502_o)
      n10976_q <= 3'b000;
    else
      n10976_q <= n9693_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1538:1  */
  assign n10977_o = {n9734_o, n10974_q, n9729_o, n10975_q, n9724_o, n10976_q};
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10978_q <= 1'b0;
    else
      n10978_q <= n10781_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10979_q <= 2'b00;
    else
      n10979_q <= n10811_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n10980_o = {n10978_q, n10859_o, n10979_q};
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10981_q <= 1'b0;
    else
      n10981_q <= n10792_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10982_q <= 2'b00;
    else
      n10982_q <= n10816_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1908:4  */
  assign n10983_o = {n10981_q, n10866_o, n10982_q};
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  assign n10984_o = n9457_o ? n9452_o : curr_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10985_q <= 1'b0;
    else
      n10985_q <= n10984_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10986_q <= 2'b00;
    else
      n10986_q <= n10460_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10987_q <= 2'b00;
    else
      n10987_q <= n10462_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1925:7  */
  always @(posedge clock_in or posedge n10356_o)
    if (n10356_o)
      n10988_q <= 1'b0;
    else
      n10988_q <= n10463_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  assign n10989_o = n9055_o ? template_r : src_template_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10990_q <= 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n10990_q <= n10989_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  assign n10991_o = load_r ? n9054_o : dest_template_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10992_q <= 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n10992_q <= n10991_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1361:9  */
  always @(posedge clock_in or posedge n9046_o)
    if (n9046_o)
      n10993_q <= 776'b00000000000000000000000011111111111111111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n10993_q <= n9458_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1352:5  */
  assign n10994_o = {n10100_o, n9991_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n10995_o = n10248_o ? task_start_addr : task_start_addr_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n10996_q <= 11'b00000000000;
    else
      n10996_q <= n10995_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n10997_o = n10248_o ? task_pcore : task_pcore_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n10998_q <= 5'b11111;
    else
      n10998_q <= n10997_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n10999_o = n10248_o ? task_tid_mask : task_tid_mask_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n11000_q <= 4'b1111;
    else
      n11000_q <= n10999_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n11001_o = n10248_o ? task_data_model : task_data_model_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n11002_q <= 2'b00;
    else
      n11002_q <= n11001_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n11003_o = n10248_o ? task_iregister_auto : task_iregister_auto_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n11004_q <= 28'b0000000000000000000000000000;
    else
      n11004_q <= n11003_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n11005_o = n10248_o ? task_lockstep : task_lockstep_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n11006_q <= 1'b0;
    else
      n11006_q <= n11005_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n11007_q <= 1'b0;
    else
      n11007_q <= n10258_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  assign n11008_o = n10248_o ? task_vm : task_vm_r;
  /* ../../HW/src/dp/dp_fetch.vhd:1835:9  */
  always @(posedge clock_in or posedge n10246_o)
    if (n10246_o)
      n11009_q <= 1'b0;
    else
      n11009_q <= n11008_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1263:7  */
  always @(posedge clock_in or posedge n8922_o)
    if (n8922_o)
      n11011_q <= 12'b000000000000;
    else
      n11011_q <= bus_waddr_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1263:7  */
  always @(posedge clock_in or posedge n8922_o)
    if (n8922_o)
      n11012_q <= 12'b000000000000;
    else
      n11012_q <= bus_raddr_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1263:7  */
  always @(posedge clock_in or posedge n8922_o)
    if (n8922_o)
      n11013_q <= 1'b0;
    else
      n11013_q <= n8926_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1263:7  */
  always @(posedge clock_in or posedge n8922_o)
    if (n8922_o)
      n11014_q <= 1'b0;
    else
      n11014_q <= bus_read_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1263:7  */
  always @(posedge clock_in or posedge n8922_o)
    if (n8922_o)
      n11015_q <= 32'b00000000000000000000000000000000;
    else
      n11015_q <= bus_writedata_in;
  /* ../../HW/src/dp/dp_fetch.vhd:1292:9  */
  always @(posedge clock_in or posedge n8947_o)
    if (n8947_o)
      n11016_q <= 1'b0;
    else
      n11016_q <= n9014_o;
  /* ../../HW/src/dp/dp_fetch.vhd:1150:20  */
  assign n11017_o = new_cmd_is_safe_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1149:20  */
  assign n11018_o = new_cmd_is_safe_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1148:21  */
  assign n11019_o = new_cmd_is_safe_r[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1147:16  */
  assign n11020_o = new_cmd_is_safe_r[3];
  /* ../../HW/src/dp/dp_fetch.vhd:1133:1  */
  assign n11021_o = new_cmd_is_safe_r[4];
  /* ../../HW/src/dp/dp_fetch.vhd:1133:1  */
  assign n11022_o = new_cmd_is_safe_r[5];
  /* ../../HW/src/dp/dp_fetch.vhd:1133:1  */
  assign n11023_o = new_cmd_is_safe_r[6];
  /* ../../HW/src/dp/dp_fetch.vhd:1133:1  */
  assign n11024_o = new_cmd_is_safe_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:1093:14  */
  assign n11025_o = new_cmd_is_safe_r[8];
  /* ../../HW/src/dp/dp_fetch.vhd:1079:1  */
  assign n11026_o = new_cmd_is_safe_r[9];
  /* ../../HW/src/dp/dp_fetch.vhd:1071:27  */
  assign n11027_o = new_cmd_is_safe_r[10];
  /* ../../HW/src/dp/dp_fetch.vhd:1070:19  */
  assign n11028_o = new_cmd_is_safe_r[11];
  /* ../../HW/src/dp/dp_fetch.vhd:1069:21  */
  assign n11029_o = new_cmd_is_safe_r[12];
  /* ../../HW/src/dp/dp_fetch.vhd:1068:21  */
  assign n11030_o = new_cmd_is_safe_r[13];
  /* ../../HW/src/dp/dp_fetch.vhd:1065:24  */
  assign n11031_o = new_cmd_is_safe_r[14];
  /* ../../HW/src/dp/dp_fetch.vhd:1064:24  */
  assign n11032_o = new_cmd_is_safe_r[15];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11033_o = {n9971_o, n9975_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11034_o = n11033_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11034_o)
      2'b00: n11035_o = n11017_o;
      2'b01: n11035_o = n11018_o;
      2'b10: n11035_o = n11019_o;
      2'b11: n11035_o = n11020_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11036_o = n11033_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11036_o)
      2'b00: n11037_o = n11021_o;
      2'b01: n11037_o = n11022_o;
      2'b10: n11037_o = n11023_o;
      2'b11: n11037_o = n11024_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11038_o = n11033_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11038_o)
      2'b00: n11039_o = n11025_o;
      2'b01: n11039_o = n11026_o;
      2'b10: n11039_o = n11027_o;
      2'b11: n11039_o = n11028_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11040_o = n11033_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11040_o)
      2'b00: n11041_o = n11029_o;
      2'b01: n11041_o = n11030_o;
      2'b10: n11041_o = n11031_o;
      2'b11: n11041_o = n11032_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11042_o = n11033_o[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11042_o)
      2'b00: n11043_o = n11035_o;
      2'b01: n11043_o = n11037_o;
      2'b10: n11043_o = n11039_o;
      2'b11: n11043_o = n11041_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11044_o = new_cmd_is_safe_r[0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:84  */
  assign n11045_o = new_cmd_is_safe_r[1];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:48  */
  assign n11046_o = new_cmd_is_safe_r[2];
  /* ../../HW/src/dp/dp_fetch.vhd:1026:1  */
  assign n11047_o = new_cmd_is_safe_r[3];
  /* ../../HW/src/dp/dp_fetch.vhd:1026:1  */
  assign n11048_o = new_cmd_is_safe_r[4];
  /* ../../HW/src/dp/dp_fetch.vhd:86:20  */
  assign n11049_o = new_cmd_is_safe_r[5];
  /* ../../HW/src/dp/dp_fetch.vhd:80:20  */
  assign n11050_o = new_cmd_is_safe_r[6];
  /* ../../HW/src/dp/dp_fetch.vhd:79:20  */
  assign n11051_o = new_cmd_is_safe_r[7];
  /* ../../HW/src/dp/dp_fetch.vhd:78:20  */
  assign n11052_o = new_cmd_is_safe_r[8];
  /* ../../HW/src/dp/dp_fetch.vhd:77:20  */
  assign n11053_o = new_cmd_is_safe_r[9];
  /* ../../HW/src/dp/dp_fetch.vhd:76:20  */
  assign n11054_o = new_cmd_is_safe_r[10];
  /* ../../HW/src/dp/dp_fetch.vhd:75:20  */
  assign n11055_o = new_cmd_is_safe_r[11];
  /* ../../HW/src/dp/dp_fetch.vhd:74:20  */
  assign n11056_o = new_cmd_is_safe_r[12];
  /* ../../HW/src/dp/dp_fetch.vhd:73:20  */
  assign n11057_o = new_cmd_is_safe_r[13];
  /* ../../HW/src/dp/dp_fetch.vhd:72:20  */
  assign n11058_o = new_cmd_is_safe_r[14];
  /* ../../HW/src/dp/dp_fetch.vhd:62:20  */
  assign n11059_o = new_cmd_is_safe_r[15];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11060_o = {n10080_o, n10084_o};
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11061_o = n11060_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11061_o)
      2'b00: n11062_o = n11044_o;
      2'b01: n11062_o = n11045_o;
      2'b10: n11062_o = n11046_o;
      2'b11: n11062_o = n11047_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11063_o = n11060_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11063_o)
      2'b00: n11064_o = n11048_o;
      2'b01: n11064_o = n11049_o;
      2'b10: n11064_o = n11050_o;
      2'b11: n11064_o = n11051_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11065_o = n11060_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11065_o)
      2'b00: n11066_o = n11052_o;
      2'b01: n11066_o = n11053_o;
      2'b10: n11066_o = n11054_o;
      2'b11: n11066_o = n11055_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11067_o = n11060_o[1:0];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11067_o)
      2'b00: n11068_o = n11056_o;
      2'b01: n11068_o = n11057_o;
      2'b10: n11068_o = n11058_o;
      2'b11: n11068_o = n11059_o;
    endcase
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  assign n11069_o = n11060_o[3:2];
  /* ../../HW/src/dp/dp_fetch.vhd:1678:83  */
  always @*
    case (n11069_o)
      2'b00: n11070_o = n11062_o;
      2'b01: n11070_o = n11064_o;
      2'b10: n11070_o = n11066_o;
      2'b11: n11070_o = n11068_o;
    endcase
endmodule

module dpram_64_64_6_6_35_35
  (input  [5:0] address_a,
   input  clock,
   input  [34:0] data_a,
   input  wren_a,
   input  [5:0] address_b,
   output [34:0] q_b);
  wire [5:0] address_r;
  reg [5:0] n7767_q;
  wire [34:0] n7768_data; // mem_rd
  assign q_b = n7768_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n7767_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n7767_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [34:0] ram_block[63:0] ; // memory
  assign n7768_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module dpram_16_16_4_4_37_37
  (input  [3:0] address_a,
   input  clock,
   input  [36:0] data_a,
   input  wren_a,
   input  [3:0] address_b,
   output [36:0] q_b);
  wire [3:0] address_r;
  reg [3:0] n7744_q;
  wire [36:0] n7745_data; // mem_rd
  assign q_b = n7745_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n7744_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n7744_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [36:0] ram_block[15:0] ; // memory
  assign n7745_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module dpram_512_512_9_9_64_64
  (input  [8:0] address_a,
   input  clock,
   input  [63:0] data_a,
   input  wren_a,
   input  [8:0] address_b,
   output [63:0] q_b);
  wire [8:0] address_r;
  reg [8:0] n7721_q;
  wire [63:0] n7722_data; // mem_rd
  assign q_b = n7722_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n7721_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n7721_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [63:0] ram_block[511:0] ; // memory
  assign n7722_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module dpram_be_2048_2048_11_11_64_64
  (input  [10:0] address_a,
   input  [7:0] byteena_a,
   input  clock0,
   input  [63:0] data_a,
   input  wren_a,
   input  [10:0] address_b,
   output [63:0] q_b);
  wire [63:0] q;
  wire [63:0] data;
  wire [10:0] address_r;
  wire [7:0] n7577_o;
  wire [7:0] n7578_o;
  wire [7:0] n7579_o;
  wire [7:0] n7580_o;
  wire [7:0] n7581_o;
  wire [7:0] n7582_o;
  wire [7:0] n7583_o;
  wire [7:0] n7584_o;
  wire [7:0] n7585_o;
  wire [7:0] n7586_o;
  wire [7:0] n7587_o;
  wire [7:0] n7588_o;
  wire [7:0] n7589_o;
  wire [7:0] n7590_o;
  wire [7:0] n7591_o;
  wire [7:0] n7592_o;
  wire n7596_o;
  wire [7:0] n7601_o;
  wire n7604_o;
  wire [7:0] n7609_o;
  wire n7612_o;
  wire [7:0] n7617_o;
  wire n7620_o;
  wire [7:0] n7625_o;
  wire n7628_o;
  wire [7:0] n7633_o;
  wire n7636_o;
  wire [7:0] n7641_o;
  wire n7644_o;
  wire [7:0] n7649_o;
  wire n7652_o;
  wire [7:0] n7657_o;
  wire n7664_o;
  wire n7666_o;
  wire n7668_o;
  wire n7670_o;
  wire n7672_o;
  wire n7674_o;
  wire n7676_o;
  wire n7678_o;
  wire [63:0] n7681_o;
  reg [10:0] n7682_q;
  wire [63:0] n7683_o;
  wire [7:0] n7684_data; // mem_rd
  wire [7:0] n7685_data; // mem_rd
  wire [7:0] n7686_data; // mem_rd
  wire [7:0] n7687_data; // mem_rd
  wire [7:0] n7688_data; // mem_rd
  wire [7:0] n7689_data; // mem_rd
  wire [7:0] n7690_data; // mem_rd
  wire [7:0] n7691_data; // mem_rd
  wire [63:0] n7692_o;
  assign q_b = n7683_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:55:8  */
  assign q = n7692_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:56:8  */
  assign data = n7681_o; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:57:8  */
  assign address_r = n7682_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7577_o = q[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7578_o = q[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7579_o = q[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7580_o = q[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7581_o = q[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7582_o = q[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7583_o = q[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:66:30  */
  assign n7584_o = q[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7585_o = data_a[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7586_o = data_a[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7587_o = data_a[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7588_o = data_a[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7589_o = data_a[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7590_o = data_a[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7591_o = data_a[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:70:21  */
  assign n7592_o = data_a[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7596_o = byteena_a[0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7601_o = data[63:56];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7604_o = byteena_a[1];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7609_o = data[55:48];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7612_o = byteena_a[2];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7617_o = data[47:40];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7620_o = byteena_a[3];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7625_o = data[39:32];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7628_o = byteena_a[4];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7633_o = data[31:24];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7636_o = byteena_a[5];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7641_o = data[23:16];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7644_o = byteena_a[6];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7649_o = data[15:8];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:78:25  */
  assign n7652_o = byteena_a[7];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:69  */
  assign n7657_o = data[7:0];
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7664_o = wren_a & n7652_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7666_o = wren_a & n7644_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7668_o = wren_a & n7636_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7670_o = wren_a & n7628_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7672_o = wren_a & n7620_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7674_o = wren_a & n7612_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7676_o = wren_a & n7604_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:30:8  */
  assign n7678_o = wren_a & n7596_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n7681_o = {n7585_o, n7586_o, n7587_o, n7588_o, n7589_o, n7590_o, n7591_o, n7592_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  always @(posedge clock0)
    n7682_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:75:4  */
  assign n7683_o = {n7584_o, n7583_o, n7582_o, n7581_o, n7580_o, n7579_o, n7578_o, n7577_o};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n1[2047:0] ; // memory
  assign n7684_data = ram_block_n1[address_r];
  always @(posedge clock0)
    if (n7664_o)
      ram_block_n1[address_a] <= n7657_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  reg [7:0] ram_block_n2[2047:0] ; // memory
  assign n7685_data = ram_block_n2[address_r];
  always @(posedge clock0)
    if (n7666_o)
      ram_block_n2[address_a] <= n7649_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n3[2047:0] ; // memory
  assign n7686_data = ram_block_n3[address_r];
  always @(posedge clock0)
    if (n7668_o)
      ram_block_n3[address_a] <= n7641_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n4[2047:0] ; // memory
  assign n7687_data = ram_block_n4[address_r];
  always @(posedge clock0)
    if (n7670_o)
      ram_block_n4[address_a] <= n7633_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n5[2047:0] ; // memory
  assign n7688_data = ram_block_n5[address_r];
  always @(posedge clock0)
    if (n7672_o)
      ram_block_n5[address_a] <= n7625_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n6[2047:0] ; // memory
  assign n7689_data = ram_block_n6[address_r];
  always @(posedge clock0)
    if (n7674_o)
      ram_block_n6[address_a] <= n7617_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n7[2047:0] ; // memory
  assign n7690_data = ram_block_n7[address_r];
  always @(posedge clock0)
    if (n7676_o)
      ram_block_n7[address_a] <= n7609_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  reg [7:0] ram_block_n8[2047:0] ; // memory
  assign n7691_data = ram_block_n8[address_r];
  always @(posedge clock0)
    if (n7678_o)
      ram_block_n8[address_a] <= n7601_o;
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:63:16  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  assign n7692_o = {n7691_data, n7690_data, n7689_data, n7688_data, n7687_data, n7686_data, n7685_data, n7684_data};
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
  /* ../../HW/platform/simulation/DPRAM_BE.vhd:79:26  */
endmodule

module delay_3
  (input  clock_in,
   input  reset_in,
   input  in_in,
   input  enable_in,
   output out_out);
  wire [2:0] fifo_r;
  wire n7549_o;
  wire n7552_o;
  wire n7557_o;
  wire n7558_o;
  wire n7559_o;
  wire n7560_o;
  wire n7561_o;
  wire n7562_o;
  wire n7563_o;
  wire n7564_o;
  wire [2:0] n7565_o;
  wire [2:0] n7567_o;
  reg [2:0] n7570_q;
  assign out_out = n7549_o;
  /* ../../HW/src/util/delay.vhd:46:8  */
  assign fifo_r = n7570_q; // (signal)
  /* ../../HW/src/util/delay.vhd:48:18  */
  assign n7549_o = fifo_r[0];
  /* ../../HW/src/util/delay.vhd:51:16  */
  assign n7552_o = ~reset_in;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n7557_o = fifo_r[1];
  /* ../../HW/platform/simulation/DPRAM.vhd:58:1  */
  assign n7558_o = fifo_r[0];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n7559_o = enable_in ? n7557_o : n7558_o;
  /* ../../HW/src/util/delay.vhd:60:44  */
  assign n7560_o = fifo_r[2];
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign n7561_o = fifo_r[1];
  /* ../../HW/src/util/delay.vhd:59:21  */
  assign n7562_o = enable_in ? n7560_o : n7561_o;
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign n7563_o = fifo_r[2];
  /* ../../HW/src/util/delay.vhd:64:13  */
  assign n7564_o = enable_in ? in_in : n7563_o;
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign n7565_o = {n7564_o, n7562_o, n7559_o};
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign n7567_o = {1'b0, 1'b0, 1'b0};
  /* ../../HW/src/util/delay.vhd:56:9  */
  always @(posedge clock_in or posedge n7552_o)
    if (n7552_o)
      n7570_q <= n7567_o;
    else
      n7570_q <= n7565_o;
endmodule

module dpram_64_64_6_6_32_32
  (input  [5:0] address_a,
   input  clock,
   input  [31:0] data_a,
   input  wren_a,
   input  [5:0] address_b,
   output [31:0] q_b);
  wire [5:0] address_r;
  reg [5:0] n7545_q;
  wire [31:0] n7546_data; // mem_rd
  assign q_b = n7546_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n7545_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n7545_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [31:0] ram_block[63:0] ; // memory
  assign n7546_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module dpram_64_64_6_6_24_24
  (input  [5:0] address_a,
   input  clock,
   input  [23:0] data_a,
   input  wren_a,
   input  [5:0] address_b,
   output [23:0] q_b);
  wire [5:0] address_r;
  reg [5:0] n7522_q;
  wire [23:0] n7523_data; // mem_rd
  assign q_b = n7523_data;
  /* ../../HW/platform/simulation/DPRAM.vhd:52:8  */
  assign address_r = n7522_q; // (signal)
  /* ../../HW/platform/simulation/DPRAM.vhd:60:4  */
  always @(posedge clock)
    n7522_q <= address_b;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  reg [23:0] ram_block[63:0] ; // memory
  assign n7523_data = ram_block[address_r];
  always @(posedge clock)
    if (wren_a)
      ram_block[address_a] <= data_a;
  /* ../../HW/platform/simulation/DPRAM.vhd:56:18  */
  /* ../../HW/platform/simulation/DPRAM.vhd:62:20  */
endmodule

module cell_1
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_fork_in,
   input  dp_rd_share_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  [3:0] enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_readdata_valid_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out,
   output [3:0] i_y_neg_out,
   output [3:0] i_y_zero_out);
  wire [3:0] dp_readena;
  wire [7:0] dp_read_data_flow;
  wire [3:0] dp_read_stream;
  wire [7:0] dp_read_stream_id;
  wire [7:0] dp_read_data_type;
  wire [3:0] dp_read_gen_valid;
  wire [95:0] dp_readdata;
  wire dp_readdata_vm;
  wire dp_readena_r;
  wire [95:0] dp_readdata_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [2:0] dp_read_vector;
  wire [2:0] dp_read_vector_r;
  wire [2:0] dp_read_vaddr;
  wire [2:0] dp_read_vaddr_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire [21:0] dp_rd_addr_step_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire [21:0] dp_wr_addr_step_in_r;
  wire dp_wr_fork_in_r;
  wire dp_wr_share_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_read_in_r;
  wire dp_rd_fork_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n7091_o;
  wire n7094_o;
  wire n7097_o;
  wire [3:0] n7098_o;
  wire n7100_o;
  wire n7103_o;
  wire [1:0] n7104_o;
  wire [1:0] n7106_o;
  wire [1:0] n7108_o;
  wire [1:0] n7109_o;
  wire [1:0] n7110_o;
  wire [1:0] n7111_o;
  wire [1:0] n7112_o;
  wire [1:0] n7113_o;
  wire n7114_o;
  wire n7116_o;
  wire n7118_o;
  wire n7119_o;
  wire n7120_o;
  wire n7121_o;
  wire n7122_o;
  wire n7123_o;
  wire [1:0] n7124_o;
  wire [1:0] n7126_o;
  wire [1:0] n7128_o;
  wire [1:0] n7129_o;
  wire [1:0] n7130_o;
  wire [1:0] n7131_o;
  wire [1:0] n7132_o;
  wire [1:0] n7133_o;
  wire [1:0] n7134_o;
  wire [1:0] n7136_o;
  wire [1:0] n7138_o;
  wire [1:0] n7139_o;
  wire [1:0] n7140_o;
  wire [1:0] n7141_o;
  wire [1:0] n7142_o;
  wire [1:0] n7143_o;
  wire n7206_o;
  wire gen_reg_n1_gen1_pcore_i_n7207;
  wire gen_reg_n1_gen1_pcore_i_n7208;
  wire [95:0] gen_reg_n1_gen1_pcore_i_n7209;
  wire gen_reg_n1_gen1_pcore_i_n7210;
  wire gen_reg_n1_gen1_pcore_i_n7211;
  wire [2:0] gen_reg_n1_gen1_pcore_i_n7212;
  wire [2:0] gen_reg_n1_gen1_pcore_i_n7213;
  wire gen_reg_n1_gen1_pcore_i_n7214;
  wire [1:0] gen_reg_n1_gen1_pcore_i_n7215;
  wire [1:0] gen_reg_n1_gen1_pcore_i_n7216;
  wire gen_reg_n1_gen1_pcore_i_n7217;
  wire [1:0] gen_reg_n1_gen1_pcore_i_n7218;
  wire gen_reg_n1_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n1_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n1_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n1_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n1_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n1_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n1_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n1_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n1_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n1_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n1_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n1_gen1_pcore_i_dp_read_stream_id_out;
  wire n7243_o;
  wire gen_reg_n2_gen1_pcore_i_n7244;
  wire gen_reg_n2_gen1_pcore_i_n7245;
  wire [95:0] gen_reg_n2_gen1_pcore_i_n7246;
  wire gen_reg_n2_gen1_pcore_i_n7247;
  wire gen_reg_n2_gen1_pcore_i_n7248;
  wire [2:0] gen_reg_n2_gen1_pcore_i_n7249;
  wire [2:0] gen_reg_n2_gen1_pcore_i_n7250;
  wire gen_reg_n2_gen1_pcore_i_n7251;
  wire [1:0] gen_reg_n2_gen1_pcore_i_n7252;
  wire [1:0] gen_reg_n2_gen1_pcore_i_n7253;
  wire gen_reg_n2_gen1_pcore_i_n7254;
  wire [1:0] gen_reg_n2_gen1_pcore_i_n7255;
  wire gen_reg_n2_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n2_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n2_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n2_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n2_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n2_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n2_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n2_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n2_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n2_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n2_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n2_gen1_pcore_i_dp_read_stream_id_out;
  wire n7280_o;
  wire gen_reg_n3_gen1_pcore_i_n7281;
  wire gen_reg_n3_gen1_pcore_i_n7282;
  wire [95:0] gen_reg_n3_gen1_pcore_i_n7283;
  wire gen_reg_n3_gen1_pcore_i_n7284;
  wire gen_reg_n3_gen1_pcore_i_n7285;
  wire [2:0] gen_reg_n3_gen1_pcore_i_n7286;
  wire [2:0] gen_reg_n3_gen1_pcore_i_n7287;
  wire gen_reg_n3_gen1_pcore_i_n7288;
  wire [1:0] gen_reg_n3_gen1_pcore_i_n7289;
  wire [1:0] gen_reg_n3_gen1_pcore_i_n7290;
  wire gen_reg_n3_gen1_pcore_i_n7291;
  wire [1:0] gen_reg_n3_gen1_pcore_i_n7292;
  wire gen_reg_n3_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n3_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n3_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n3_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n3_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n3_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n3_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n3_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n3_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n3_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n3_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n3_gen1_pcore_i_dp_read_stream_id_out;
  wire n7317_o;
  wire gen_reg_n4_gen1_pcore_i_n7318;
  wire gen_reg_n4_gen1_pcore_i_n7319;
  wire [95:0] gen_reg_n4_gen1_pcore_i_n7320;
  wire gen_reg_n4_gen1_pcore_i_n7321;
  wire gen_reg_n4_gen1_pcore_i_n7322;
  wire [2:0] gen_reg_n4_gen1_pcore_i_n7323;
  wire [2:0] gen_reg_n4_gen1_pcore_i_n7324;
  wire gen_reg_n4_gen1_pcore_i_n7325;
  wire [1:0] gen_reg_n4_gen1_pcore_i_n7326;
  wire [1:0] gen_reg_n4_gen1_pcore_i_n7327;
  wire gen_reg_n4_gen1_pcore_i_n7328;
  wire [1:0] gen_reg_n4_gen1_pcore_i_n7329;
  wire gen_reg_n4_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n4_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n4_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n4_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n4_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n4_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n4_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n4_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n4_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n4_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n4_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n4_gen1_pcore_i_dp_read_stream_id_out;
  wire n7356_o;
  wire [3:0] n7437_o;
  wire [7:0] n7438_o;
  wire [3:0] n7439_o;
  wire [7:0] n7440_o;
  wire [7:0] n7441_o;
  wire [3:0] n7442_o;
  wire [95:0] n7443_o;
  wire [95:0] n7444_o;
  wire [95:0] n7445_o;
  wire n7446_o;
  wire n7447_o;
  wire n7448_o;
  reg n7449_q;
  reg [95:0] n7450_q;
  reg n7451_q;
  reg n7452_q;
  reg [1:0] n7453_q;
  reg [1:0] n7454_q;
  reg n7455_q;
  reg [1:0] n7456_q;
  wire [2:0] n7457_o;
  wire [2:0] n7458_o;
  wire [2:0] n7459_o;
  reg [2:0] n7460_q;
  wire [2:0] n7461_o;
  wire [2:0] n7462_o;
  wire [2:0] n7463_o;
  reg [2:0] n7464_q;
  reg n7465_q;
  reg n7466_q;
  reg n7467_q;
  reg [21:0] n7468_q;
  reg [21:0] n7469_q;
  reg n7470_q;
  reg [21:0] n7471_q;
  reg [21:0] n7472_q;
  reg n7473_q;
  reg n7474_q;
  reg [5:0] n7475_q;
  reg n7476_q;
  reg n7477_q;
  reg [2:0] n7478_q;
  reg [1:0] n7479_q;
  reg n7480_q;
  reg n7481_q;
  reg [2:0] n7482_q;
  reg [1:0] n7483_q;
  reg n7484_q;
  reg [1:0] n7485_q;
  reg [1:0] n7486_q;
  reg n7487_q;
  reg [1:0] n7488_q;
  reg [95:0] n7489_q;
  reg n7490_q;
  wire [95:0] n7491_o;
  wire n7492_o;
  wire [2:0] n7493_o;
  wire [2:0] n7494_o;
  wire n7495_o;
  wire [1:0] n7496_o;
  wire [1:0] n7497_o;
  wire n7498_o;
  wire [1:0] n7499_o;
  wire [3:0] n7500_o;
  wire [3:0] n7501_o;
  assign dp_readdata_out = n7491_o;
  assign dp_readdata_vm_out = n7492_o;
  assign dp_read_vector_out = n7493_o;
  assign dp_read_vaddr_out = n7494_o;
  assign dp_readdata_valid_out = dp_readena_r;
  assign dp_read_gen_valid_out = n7495_o;
  assign dp_read_data_flow_out = n7496_o;
  assign dp_read_data_type_out = n7497_o;
  assign dp_read_stream_out = n7498_o;
  assign dp_read_stream_id_out = n7499_o;
  assign i_y_neg_out = n7500_o;
  assign i_y_zero_out = n7501_o;
  /* ../../HW/src/top/cell.vhd:101:8  */
  assign dp_readena = n7437_o; // (signal)
  /* ../../HW/src/top/cell.vhd:102:8  */
  assign dp_read_data_flow = n7438_o; // (signal)
  /* ../../HW/src/top/cell.vhd:103:8  */
  assign dp_read_stream = n7439_o; // (signal)
  /* ../../HW/src/top/cell.vhd:104:8  */
  assign dp_read_stream_id = n7440_o; // (signal)
  /* ../../HW/src/top/cell.vhd:105:8  */
  assign dp_read_data_type = n7441_o; // (signal)
  /* ../../HW/src/top/cell.vhd:106:8  */
  assign dp_read_gen_valid = n7442_o; // (signal)
  /* ../../HW/src/top/cell.vhd:107:8  */
  assign dp_readdata = n7445_o; // (signal)
  /* ../../HW/src/top/cell.vhd:108:8  */
  assign dp_readdata_vm = n7448_o; // (signal)
  /* ../../HW/src/top/cell.vhd:109:8  */
  assign dp_readena_r = n7449_q; // (signal)
  /* ../../HW/src/top/cell.vhd:110:8  */
  assign dp_readdata_r = n7450_q; // (signal)
  /* ../../HW/src/top/cell.vhd:111:8  */
  assign dp_readdata_vm_r = n7451_q; // (signal)
  /* ../../HW/src/top/cell.vhd:112:8  */
  assign dp_read_gen_valid_r = n7452_q; // (signal)
  /* ../../HW/src/top/cell.vhd:113:8  */
  assign dp_read_data_flow_r = n7453_q; // (signal)
  /* ../../HW/src/top/cell.vhd:114:8  */
  assign dp_read_data_type_r = n7454_q; // (signal)
  /* ../../HW/src/top/cell.vhd:115:8  */
  assign dp_read_stream_r = n7455_q; // (signal)
  /* ../../HW/src/top/cell.vhd:116:8  */
  assign dp_read_stream_id_r = n7456_q; // (signal)
  /* ../../HW/src/top/cell.vhd:117:8  */
  assign dp_read_vector = n7459_o; // (signal)
  /* ../../HW/src/top/cell.vhd:118:8  */
  assign dp_read_vector_r = n7460_q; // (signal)
  /* ../../HW/src/top/cell.vhd:119:8  */
  assign dp_read_vaddr = n7463_o; // (signal)
  /* ../../HW/src/top/cell.vhd:120:8  */
  assign dp_read_vaddr_r = n7464_q; // (signal)
  /* ../../HW/src/top/cell.vhd:122:8  */
  assign dp_rd_vm_in_r = n7465_q; // (signal)
  /* ../../HW/src/top/cell.vhd:123:8  */
  assign dp_wr_vm_in_r = n7466_q; // (signal)
  /* ../../HW/src/top/cell.vhd:124:8  */
  assign dp_code_in_r = n7467_q; // (signal)
  /* ../../HW/src/top/cell.vhd:125:8  */
  assign dp_rd_addr_in_r = n7468_q; // (signal)
  /* ../../HW/src/top/cell.vhd:126:8  */
  assign dp_rd_addr_step_in_r = n7469_q; // (signal)
  /* ../../HW/src/top/cell.vhd:127:8  */
  assign dp_rd_share_in_r = n7470_q; // (signal)
  /* ../../HW/src/top/cell.vhd:128:8  */
  assign dp_wr_addr_in_r = n7471_q; // (signal)
  /* ../../HW/src/top/cell.vhd:129:8  */
  assign dp_wr_addr_step_in_r = n7472_q; // (signal)
  /* ../../HW/src/top/cell.vhd:130:8  */
  assign dp_wr_fork_in_r = n7473_q; // (signal)
  /* ../../HW/src/top/cell.vhd:131:8  */
  assign dp_wr_share_in_r = n7474_q; // (signal)
  /* ../../HW/src/top/cell.vhd:132:8  */
  assign dp_wr_mcast_in_r = n7475_q; // (signal)
  /* ../../HW/src/top/cell.vhd:133:8  */
  assign dp_write_in_r = n7476_q; // (signal)
  /* ../../HW/src/top/cell.vhd:134:8  */
  assign dp_write_gen_valid_in_r = n7477_q; // (signal)
  /* ../../HW/src/top/cell.vhd:135:8  */
  assign dp_write_vector_in_r = n7478_q; // (signal)
  /* ../../HW/src/top/cell.vhd:136:8  */
  assign dp_write_scatter_in_r = n7479_q; // (signal)
  /* ../../HW/src/top/cell.vhd:137:8  */
  assign dp_read_in_r = n7480_q; // (signal)
  /* ../../HW/src/top/cell.vhd:138:8  */
  assign dp_rd_fork_in_r = n7481_q; // (signal)
  /* ../../HW/src/top/cell.vhd:139:8  */
  assign dp_read_vector_in_r = n7482_q; // (signal)
  /* ../../HW/src/top/cell.vhd:140:8  */
  assign dp_read_scatter_in_r = n7483_q; // (signal)
  /* ../../HW/src/top/cell.vhd:141:8  */
  assign dp_read_gen_valid_in_r = n7484_q; // (signal)
  /* ../../HW/src/top/cell.vhd:142:8  */
  assign dp_read_data_flow_in_r = n7485_q; // (signal)
  /* ../../HW/src/top/cell.vhd:143:8  */
  assign dp_read_data_type_in_r = n7486_q; // (signal)
  /* ../../HW/src/top/cell.vhd:144:8  */
  assign dp_read_stream_in_r = n7487_q; // (signal)
  /* ../../HW/src/top/cell.vhd:145:8  */
  assign dp_read_stream_id_in_r = n7488_q; // (signal)
  /* ../../HW/src/top/cell.vhd:146:8  */
  assign dp_writedata_in_r = n7489_q; // (signal)
  /* ../../HW/src/top/cell.vhd:147:8  */
  assign dp_config_in_r = n7490_q; // (signal)
  /* ../../HW/src/top/cell.vhd:170:16  */
  assign n7091_o = ~reset_in;
  /* ../../HW/src/top/cell.vhd:184:27  */
  assign n7094_o = dp_readena == 4'b0000;
  /* ../../HW/src/top/cell.vhd:184:13  */
  assign n7097_o = n7094_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/cell.vhd:189:48  */
  assign n7098_o = dp_readena & dp_read_gen_valid;
  /* ../../HW/src/top/cell.vhd:190:36  */
  assign n7100_o = n7098_o == 4'b0000;
  /* ../../HW/src/top/cell.vhd:190:13  */
  assign n7103_o = n7100_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n7104_o = dp_read_data_flow[1:0];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n7106_o = 2'b00 | n7104_o;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n7108_o = dp_read_data_flow[3:2];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n7109_o = n7106_o | n7108_o;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n7110_o = dp_read_data_flow[5:4];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n7111_o = n7109_o | n7110_o;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n7112_o = dp_read_data_flow[7:6];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n7113_o = n7111_o | n7112_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n7114_o = dp_read_stream[0];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n7116_o = 1'b0 | n7114_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n7118_o = dp_read_stream[1];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n7119_o = n7116_o | n7118_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n7120_o = dp_read_stream[2];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n7121_o = n7119_o | n7120_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n7122_o = dp_read_stream[3];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n7123_o = n7121_o | n7122_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n7124_o = dp_read_stream_id[1:0];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n7126_o = 2'b00 | n7124_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n7128_o = dp_read_stream_id[3:2];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n7129_o = n7126_o | n7128_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n7130_o = dp_read_stream_id[5:4];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n7131_o = n7129_o | n7130_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n7132_o = dp_read_stream_id[7:6];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n7133_o = n7131_o | n7132_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n7134_o = dp_read_data_type[1:0];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n7136_o = 2'b00 | n7134_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n7138_o = dp_read_data_type[3:2];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n7139_o = n7136_o | n7138_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n7140_o = dp_read_data_type[5:4];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n7141_o = n7139_o | n7140_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n7142_o = dp_read_data_type[7:6];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n7143_o = n7141_o | n7142_o;
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n7206_o = enable_in[0];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n1_gen1_pcore_i_n7207 = gen_reg_n1_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n1_gen1_pcore_i_n7208 = gen_reg_n1_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n1_gen1_pcore_i_n7209 = gen_reg_n1_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n1_gen1_pcore_i_n7210 = gen_reg_n1_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n1_gen1_pcore_i_n7211 = gen_reg_n1_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n1_gen1_pcore_i_n7212 = gen_reg_n1_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n1_gen1_pcore_i_n7213 = gen_reg_n1_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n1_gen1_pcore_i_n7214 = gen_reg_n1_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n1_gen1_pcore_i_n7215 = gen_reg_n1_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n1_gen1_pcore_i_n7216 = gen_reg_n1_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n1_gen1_pcore_i_n7217 = gen_reg_n1_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n1_gen1_pcore_i_n7218 = gen_reg_n1_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_1_0 gen_reg_n1_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n7206_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n1_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n1_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n1_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n1_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n1_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n1_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n1_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n1_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n1_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n1_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n1_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n1_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n7243_o = enable_in[1];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n2_gen1_pcore_i_n7244 = gen_reg_n2_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n2_gen1_pcore_i_n7245 = gen_reg_n2_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n2_gen1_pcore_i_n7246 = gen_reg_n2_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n2_gen1_pcore_i_n7247 = gen_reg_n2_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n2_gen1_pcore_i_n7248 = gen_reg_n2_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n2_gen1_pcore_i_n7249 = gen_reg_n2_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n2_gen1_pcore_i_n7250 = gen_reg_n2_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n2_gen1_pcore_i_n7251 = gen_reg_n2_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n2_gen1_pcore_i_n7252 = gen_reg_n2_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n2_gen1_pcore_i_n7253 = gen_reg_n2_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n2_gen1_pcore_i_n7254 = gen_reg_n2_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n2_gen1_pcore_i_n7255 = gen_reg_n2_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_1_1 gen_reg_n2_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n7243_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n2_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n2_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n2_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n2_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n2_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n2_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n2_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n2_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n2_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n2_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n2_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n2_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n7280_o = enable_in[2];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n3_gen1_pcore_i_n7281 = gen_reg_n3_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n3_gen1_pcore_i_n7282 = gen_reg_n3_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n3_gen1_pcore_i_n7283 = gen_reg_n3_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n3_gen1_pcore_i_n7284 = gen_reg_n3_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n3_gen1_pcore_i_n7285 = gen_reg_n3_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n3_gen1_pcore_i_n7286 = gen_reg_n3_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n3_gen1_pcore_i_n7287 = gen_reg_n3_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n3_gen1_pcore_i_n7288 = gen_reg_n3_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n3_gen1_pcore_i_n7289 = gen_reg_n3_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n3_gen1_pcore_i_n7290 = gen_reg_n3_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n3_gen1_pcore_i_n7291 = gen_reg_n3_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n3_gen1_pcore_i_n7292 = gen_reg_n3_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_1_2 gen_reg_n3_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n7280_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n3_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n3_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n3_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n3_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n3_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n3_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n3_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n3_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n3_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n3_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n3_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n3_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n7317_o = enable_in[3];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n4_gen1_pcore_i_n7318 = gen_reg_n4_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n4_gen1_pcore_i_n7319 = gen_reg_n4_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n4_gen1_pcore_i_n7320 = gen_reg_n4_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n4_gen1_pcore_i_n7321 = gen_reg_n4_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n4_gen1_pcore_i_n7322 = gen_reg_n4_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n4_gen1_pcore_i_n7323 = gen_reg_n4_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n4_gen1_pcore_i_n7324 = gen_reg_n4_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n4_gen1_pcore_i_n7325 = gen_reg_n4_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n4_gen1_pcore_i_n7326 = gen_reg_n4_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n4_gen1_pcore_i_n7327 = gen_reg_n4_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n4_gen1_pcore_i_n7328 = gen_reg_n4_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n4_gen1_pcore_i_n7329 = gen_reg_n4_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_1_3 gen_reg_n4_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n7317_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n4_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n4_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n4_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n4_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n4_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n4_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n4_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n4_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n4_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n4_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n4_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n4_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:322:13  */
  assign n7356_o = ~reset_in;
  assign n7437_o = {gen_reg_n4_gen1_pcore_i_n7322, gen_reg_n3_gen1_pcore_i_n7285, gen_reg_n2_gen1_pcore_i_n7248, gen_reg_n1_gen1_pcore_i_n7211};
  assign n7438_o = {gen_reg_n4_gen1_pcore_i_n7326, gen_reg_n3_gen1_pcore_i_n7289, gen_reg_n2_gen1_pcore_i_n7252, gen_reg_n1_gen1_pcore_i_n7215};
  assign n7439_o = {gen_reg_n4_gen1_pcore_i_n7328, gen_reg_n3_gen1_pcore_i_n7291, gen_reg_n2_gen1_pcore_i_n7254, gen_reg_n1_gen1_pcore_i_n7217};
  assign n7440_o = {gen_reg_n4_gen1_pcore_i_n7329, gen_reg_n3_gen1_pcore_i_n7292, gen_reg_n2_gen1_pcore_i_n7255, gen_reg_n1_gen1_pcore_i_n7218};
  assign n7441_o = {gen_reg_n4_gen1_pcore_i_n7327, gen_reg_n3_gen1_pcore_i_n7290, gen_reg_n2_gen1_pcore_i_n7253, gen_reg_n1_gen1_pcore_i_n7216};
  assign n7442_o = {gen_reg_n4_gen1_pcore_i_n7325, gen_reg_n3_gen1_pcore_i_n7288, gen_reg_n2_gen1_pcore_i_n7251, gen_reg_n1_gen1_pcore_i_n7214};
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7443_o = gen_reg_n1_gen1_pcore_i_n7209;
  assign n7443_o = gen_reg_n2_gen1_pcore_i_n7246;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7444_o = n7443_o;
  assign n7444_o = gen_reg_n3_gen1_pcore_i_n7283;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7445_o = n7444_o;
  assign n7445_o = gen_reg_n4_gen1_pcore_i_n7320;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7446_o = gen_reg_n1_gen1_pcore_i_n7210;
  assign n7446_o = gen_reg_n2_gen1_pcore_i_n7247;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7447_o = n7446_o;
  assign n7447_o = gen_reg_n3_gen1_pcore_i_n7284;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7448_o = n7447_o;
  assign n7448_o = gen_reg_n4_gen1_pcore_i_n7321;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7449_q <= 1'b0;
    else
      n7449_q <= n7097_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7450_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n7450_q <= dp_readdata;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7451_q <= 1'b0;
    else
      n7451_q <= dp_readdata_vm;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7452_q <= 1'b0;
    else
      n7452_q <= n7103_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7453_q <= 2'b00;
    else
      n7453_q <= n7113_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7454_q <= 2'b00;
    else
      n7454_q <= n7143_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7455_q <= 1'b0;
    else
      n7455_q <= n7123_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7456_q <= 2'b00;
    else
      n7456_q <= n7133_o;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7457_o = gen_reg_n1_gen1_pcore_i_n7212;
  assign n7457_o = gen_reg_n2_gen1_pcore_i_n7249;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7458_o = n7457_o;
  assign n7458_o = gen_reg_n3_gen1_pcore_i_n7286;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7459_o = n7458_o;
  assign n7459_o = gen_reg_n4_gen1_pcore_i_n7323;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7460_q <= 3'b000;
    else
      n7460_q <= dp_read_vector;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7461_o = gen_reg_n1_gen1_pcore_i_n7213;
  assign n7461_o = gen_reg_n2_gen1_pcore_i_n7250;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7462_o = n7461_o;
  assign n7462_o = gen_reg_n3_gen1_pcore_i_n7287;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7463_o = n7462_o;
  assign n7463_o = gen_reg_n4_gen1_pcore_i_n7324;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n7091_o)
    if (n7091_o)
      n7464_q <= 3'b000;
    else
      n7464_q <= dp_read_vaddr;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7465_q <= 1'b0;
    else
      n7465_q <= dp_rd_vm_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7466_q <= 1'b0;
    else
      n7466_q <= dp_wr_vm_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7467_q <= 1'b0;
    else
      n7467_q <= dp_code_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7468_q <= 22'b0000000000000000000000;
    else
      n7468_q <= dp_rd_addr_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7469_q <= 22'b0000000000000000000000;
    else
      n7469_q <= dp_rd_addr_step_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7470_q <= 1'b0;
    else
      n7470_q <= dp_rd_share_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7471_q <= 22'b0000000000000000000000;
    else
      n7471_q <= dp_wr_addr_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7472_q <= 22'b0000000000000000000000;
    else
      n7472_q <= dp_wr_addr_step_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7473_q <= 1'b0;
    else
      n7473_q <= dp_wr_fork_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7474_q <= 1'b0;
    else
      n7474_q <= dp_wr_share_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7475_q <= 6'b000000;
    else
      n7475_q <= dp_wr_mcast_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7476_q <= 1'b0;
    else
      n7476_q <= dp_write_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7477_q <= 1'b0;
    else
      n7477_q <= dp_write_gen_valid_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7478_q <= 3'b000;
    else
      n7478_q <= dp_write_vector_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7479_q <= 2'b00;
    else
      n7479_q <= dp_write_scatter_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7480_q <= 1'b0;
    else
      n7480_q <= dp_read_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7481_q <= 1'b0;
    else
      n7481_q <= dp_rd_fork_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7482_q <= 3'b000;
    else
      n7482_q <= dp_read_vector_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7483_q <= 2'b00;
    else
      n7483_q <= dp_read_scatter_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7484_q <= 1'b0;
    else
      n7484_q <= dp_read_gen_valid_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7485_q <= 2'b00;
    else
      n7485_q <= dp_read_data_flow_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7486_q <= 2'b00;
    else
      n7486_q <= dp_read_data_type_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7487_q <= 1'b0;
    else
      n7487_q <= dp_read_stream_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7488_q <= 2'b00;
    else
      n7488_q <= dp_read_stream_id_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7489_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n7489_q <= dp_writedata_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n7356_o)
    if (n7356_o)
      n7490_q <= 1'b0;
    else
      n7490_q <= dp_config_in;
  /* ../../HW/src/top/cell.vhd:151:34  */
  assign n7491_o = dp_readena_r ? dp_readdata_r : 96'bz;
  /* ../../HW/src/top/cell.vhd:152:40  */
  assign n7492_o = dp_readena_r ? dp_readdata_vm_r : 1'bz;
  /* ../../HW/src/top/cell.vhd:159:40  */
  assign n7493_o = dp_readena_r ? dp_read_vector_r : 3'bz;
  /* ../../HW/src/top/cell.vhd:160:38  */
  assign n7494_o = dp_readena_r ? dp_read_vaddr_r : 3'bz;
  /* ../../HW/src/top/cell.vhd:154:46  */
  assign n7495_o = dp_readena_r ? dp_read_gen_valid_r : 1'bz;
  /* ../../HW/src/top/cell.vhd:155:46  */
  assign n7496_o = dp_readena_r ? dp_read_data_flow_r : 2'bz;
  /* ../../HW/src/top/cell.vhd:158:46  */
  assign n7497_o = dp_readena_r ? dp_read_data_type_r : 2'bz;
  /* ../../HW/src/top/cell.vhd:156:40  */
  assign n7498_o = dp_readena_r ? dp_read_stream_r : 1'bz;
  /* ../../HW/src/top/cell.vhd:157:46  */
  assign n7499_o = dp_readena_r ? dp_read_stream_id_r : 2'bz;
  /* ../../HW/src/top/cell.vhd:157:46  */
  assign n7500_o = {gen_reg_n4_gen1_pcore_i_n7318, gen_reg_n3_gen1_pcore_i_n7281, gen_reg_n2_gen1_pcore_i_n7244, gen_reg_n1_gen1_pcore_i_n7207};
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7501_o = {gen_reg_n4_gen1_pcore_i_n7319, gen_reg_n3_gen1_pcore_i_n7282, gen_reg_n2_gen1_pcore_i_n7245, gen_reg_n1_gen1_pcore_i_n7208};
endmodule

module cell_0
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  dp_rd_vm_in,
   input  dp_wr_vm_in,
   input  dp_code_in,
   input  [21:0] dp_rd_addr_in,
   input  [21:0] dp_rd_addr_step_in,
   input  dp_rd_fork_in,
   input  dp_rd_share_in,
   input  [21:0] dp_wr_addr_in,
   input  [21:0] dp_wr_addr_step_in,
   input  dp_wr_fork_in,
   input  dp_wr_share_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  dp_read_gen_valid_in,
   input  [1:0] dp_read_data_flow_in,
   input  [1:0] dp_read_data_type_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [95:0] dp_writedata_in,
   input  dp_config_in,
   input  [79:0] instruction_mu_in,
   input  [31:0] instruction_imu_in,
   input  instruction_mu_valid_in,
   input  instruction_imu_valid_in,
   input  vm_in,
   input  [1:0] data_model_in,
   input  [3:0] enable_in,
   input  [3:0] tid_in,
   input  tid_valid1_in,
   input  [3:0] pre_tid_in,
   input  pre_tid_valid1_in,
   input  [3:0] pre_pre_tid_in,
   input  pre_pre_tid_valid1_in,
   input  pre_pre_vm_in,
   input  [1:0] pre_pre_data_model_in,
   input  [27:0] pre_iregister_auto_in,
   output [95:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output [2:0] dp_read_vector_out,
   output [2:0] dp_read_vaddr_out,
   output dp_readdata_valid_out,
   output dp_read_gen_valid_out,
   output [1:0] dp_read_data_flow_out,
   output [1:0] dp_read_data_type_out,
   output dp_read_stream_out,
   output [1:0] dp_read_stream_id_out,
   output [3:0] i_y_neg_out,
   output [3:0] i_y_zero_out);
  wire [3:0] dp_readena;
  wire [7:0] dp_read_data_flow;
  wire [3:0] dp_read_stream;
  wire [7:0] dp_read_stream_id;
  wire [7:0] dp_read_data_type;
  wire [3:0] dp_read_gen_valid;
  wire [95:0] dp_readdata;
  wire dp_readdata_vm;
  wire dp_readena_r;
  wire [95:0] dp_readdata_r;
  wire dp_readdata_vm_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [2:0] dp_read_vector;
  wire [2:0] dp_read_vector_r;
  wire [2:0] dp_read_vaddr;
  wire [2:0] dp_read_vaddr_r;
  wire dp_rd_vm_in_r;
  wire dp_wr_vm_in_r;
  wire dp_code_in_r;
  wire [21:0] dp_rd_addr_in_r;
  wire [21:0] dp_rd_addr_step_in_r;
  wire dp_rd_share_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire [21:0] dp_wr_addr_step_in_r;
  wire dp_wr_fork_in_r;
  wire dp_wr_share_in_r;
  wire [5:0] dp_wr_mcast_in_r;
  wire dp_write_in_r;
  wire dp_write_gen_valid_in_r;
  wire [2:0] dp_write_vector_in_r;
  wire [1:0] dp_write_scatter_in_r;
  wire dp_read_in_r;
  wire dp_rd_fork_in_r;
  wire [2:0] dp_read_vector_in_r;
  wire [1:0] dp_read_scatter_in_r;
  wire dp_read_gen_valid_in_r;
  wire [1:0] dp_read_data_flow_in_r;
  wire [1:0] dp_read_data_type_in_r;
  wire dp_read_stream_in_r;
  wire [1:0] dp_read_stream_id_in_r;
  wire [95:0] dp_writedata_in_r;
  wire dp_config_in_r;
  wire n6642_o;
  wire n6645_o;
  wire n6648_o;
  wire [3:0] n6649_o;
  wire n6651_o;
  wire n6654_o;
  wire [1:0] n6655_o;
  wire [1:0] n6657_o;
  wire [1:0] n6659_o;
  wire [1:0] n6660_o;
  wire [1:0] n6661_o;
  wire [1:0] n6662_o;
  wire [1:0] n6663_o;
  wire [1:0] n6664_o;
  wire n6665_o;
  wire n6667_o;
  wire n6669_o;
  wire n6670_o;
  wire n6671_o;
  wire n6672_o;
  wire n6673_o;
  wire n6674_o;
  wire [1:0] n6675_o;
  wire [1:0] n6677_o;
  wire [1:0] n6679_o;
  wire [1:0] n6680_o;
  wire [1:0] n6681_o;
  wire [1:0] n6682_o;
  wire [1:0] n6683_o;
  wire [1:0] n6684_o;
  wire [1:0] n6685_o;
  wire [1:0] n6687_o;
  wire [1:0] n6689_o;
  wire [1:0] n6690_o;
  wire [1:0] n6691_o;
  wire [1:0] n6692_o;
  wire [1:0] n6693_o;
  wire [1:0] n6694_o;
  wire n6757_o;
  wire gen_reg_n1_gen1_pcore_i_n6758;
  wire gen_reg_n1_gen1_pcore_i_n6759;
  wire [95:0] gen_reg_n1_gen1_pcore_i_n6760;
  wire gen_reg_n1_gen1_pcore_i_n6761;
  wire gen_reg_n1_gen1_pcore_i_n6762;
  wire [2:0] gen_reg_n1_gen1_pcore_i_n6763;
  wire [2:0] gen_reg_n1_gen1_pcore_i_n6764;
  wire gen_reg_n1_gen1_pcore_i_n6765;
  wire [1:0] gen_reg_n1_gen1_pcore_i_n6766;
  wire [1:0] gen_reg_n1_gen1_pcore_i_n6767;
  wire gen_reg_n1_gen1_pcore_i_n6768;
  wire [1:0] gen_reg_n1_gen1_pcore_i_n6769;
  wire gen_reg_n1_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n1_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n1_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n1_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n1_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n1_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n1_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n1_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n1_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n1_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n1_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n1_gen1_pcore_i_dp_read_stream_id_out;
  wire n6794_o;
  wire gen_reg_n2_gen1_pcore_i_n6795;
  wire gen_reg_n2_gen1_pcore_i_n6796;
  wire [95:0] gen_reg_n2_gen1_pcore_i_n6797;
  wire gen_reg_n2_gen1_pcore_i_n6798;
  wire gen_reg_n2_gen1_pcore_i_n6799;
  wire [2:0] gen_reg_n2_gen1_pcore_i_n6800;
  wire [2:0] gen_reg_n2_gen1_pcore_i_n6801;
  wire gen_reg_n2_gen1_pcore_i_n6802;
  wire [1:0] gen_reg_n2_gen1_pcore_i_n6803;
  wire [1:0] gen_reg_n2_gen1_pcore_i_n6804;
  wire gen_reg_n2_gen1_pcore_i_n6805;
  wire [1:0] gen_reg_n2_gen1_pcore_i_n6806;
  wire gen_reg_n2_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n2_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n2_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n2_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n2_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n2_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n2_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n2_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n2_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n2_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n2_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n2_gen1_pcore_i_dp_read_stream_id_out;
  wire n6831_o;
  wire gen_reg_n3_gen1_pcore_i_n6832;
  wire gen_reg_n3_gen1_pcore_i_n6833;
  wire [95:0] gen_reg_n3_gen1_pcore_i_n6834;
  wire gen_reg_n3_gen1_pcore_i_n6835;
  wire gen_reg_n3_gen1_pcore_i_n6836;
  wire [2:0] gen_reg_n3_gen1_pcore_i_n6837;
  wire [2:0] gen_reg_n3_gen1_pcore_i_n6838;
  wire gen_reg_n3_gen1_pcore_i_n6839;
  wire [1:0] gen_reg_n3_gen1_pcore_i_n6840;
  wire [1:0] gen_reg_n3_gen1_pcore_i_n6841;
  wire gen_reg_n3_gen1_pcore_i_n6842;
  wire [1:0] gen_reg_n3_gen1_pcore_i_n6843;
  wire gen_reg_n3_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n3_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n3_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n3_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n3_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n3_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n3_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n3_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n3_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n3_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n3_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n3_gen1_pcore_i_dp_read_stream_id_out;
  wire n6868_o;
  wire gen_reg_n4_gen1_pcore_i_n6869;
  wire gen_reg_n4_gen1_pcore_i_n6870;
  wire [95:0] gen_reg_n4_gen1_pcore_i_n6871;
  wire gen_reg_n4_gen1_pcore_i_n6872;
  wire gen_reg_n4_gen1_pcore_i_n6873;
  wire [2:0] gen_reg_n4_gen1_pcore_i_n6874;
  wire [2:0] gen_reg_n4_gen1_pcore_i_n6875;
  wire gen_reg_n4_gen1_pcore_i_n6876;
  wire [1:0] gen_reg_n4_gen1_pcore_i_n6877;
  wire [1:0] gen_reg_n4_gen1_pcore_i_n6878;
  wire gen_reg_n4_gen1_pcore_i_n6879;
  wire [1:0] gen_reg_n4_gen1_pcore_i_n6880;
  wire gen_reg_n4_gen1_pcore_i_i_y_neg_out;
  wire gen_reg_n4_gen1_pcore_i_i_y_zero_out;
  wire [95:0] gen_reg_n4_gen1_pcore_i_dp_readdata_out;
  wire gen_reg_n4_gen1_pcore_i_dp_readdata_vm_out;
  wire gen_reg_n4_gen1_pcore_i_dp_readena_out;
  wire [2:0] gen_reg_n4_gen1_pcore_i_dp_read_vector_out;
  wire [2:0] gen_reg_n4_gen1_pcore_i_dp_read_vaddr_out;
  wire gen_reg_n4_gen1_pcore_i_dp_read_gen_valid_out;
  wire [1:0] gen_reg_n4_gen1_pcore_i_dp_read_data_flow_out;
  wire [1:0] gen_reg_n4_gen1_pcore_i_dp_read_data_type_out;
  wire gen_reg_n4_gen1_pcore_i_dp_read_stream_out;
  wire [1:0] gen_reg_n4_gen1_pcore_i_dp_read_stream_id_out;
  wire n6907_o;
  wire [3:0] n6988_o;
  wire [7:0] n6989_o;
  wire [3:0] n6990_o;
  wire [7:0] n6991_o;
  wire [7:0] n6992_o;
  wire [3:0] n6993_o;
  wire [95:0] n6994_o;
  wire [95:0] n6995_o;
  wire [95:0] n6996_o;
  wire n6997_o;
  wire n6998_o;
  wire n6999_o;
  reg n7000_q;
  reg [95:0] n7001_q;
  reg n7002_q;
  reg n7003_q;
  reg [1:0] n7004_q;
  reg [1:0] n7005_q;
  reg n7006_q;
  reg [1:0] n7007_q;
  wire [2:0] n7008_o;
  wire [2:0] n7009_o;
  wire [2:0] n7010_o;
  reg [2:0] n7011_q;
  wire [2:0] n7012_o;
  wire [2:0] n7013_o;
  wire [2:0] n7014_o;
  reg [2:0] n7015_q;
  reg n7016_q;
  reg n7017_q;
  reg n7018_q;
  reg [21:0] n7019_q;
  reg [21:0] n7020_q;
  reg n7021_q;
  reg [21:0] n7022_q;
  reg [21:0] n7023_q;
  reg n7024_q;
  reg n7025_q;
  reg [5:0] n7026_q;
  reg n7027_q;
  reg n7028_q;
  reg [2:0] n7029_q;
  reg [1:0] n7030_q;
  reg n7031_q;
  reg n7032_q;
  reg [2:0] n7033_q;
  reg [1:0] n7034_q;
  reg n7035_q;
  reg [1:0] n7036_q;
  reg [1:0] n7037_q;
  reg n7038_q;
  reg [1:0] n7039_q;
  reg [95:0] n7040_q;
  reg n7041_q;
  wire [95:0] n7042_o;
  wire n7043_o;
  wire [2:0] n7044_o;
  wire [2:0] n7045_o;
  wire n7046_o;
  wire [1:0] n7047_o;
  wire [1:0] n7048_o;
  wire n7049_o;
  wire [1:0] n7050_o;
  wire [3:0] n7051_o;
  wire [3:0] n7052_o;
  assign dp_readdata_out = n7042_o;
  assign dp_readdata_vm_out = n7043_o;
  assign dp_read_vector_out = n7044_o;
  assign dp_read_vaddr_out = n7045_o;
  assign dp_readdata_valid_out = dp_readena_r;
  assign dp_read_gen_valid_out = n7046_o;
  assign dp_read_data_flow_out = n7047_o;
  assign dp_read_data_type_out = n7048_o;
  assign dp_read_stream_out = n7049_o;
  assign dp_read_stream_id_out = n7050_o;
  assign i_y_neg_out = n7051_o;
  assign i_y_zero_out = n7052_o;
  /* ../../HW/src/top/cell.vhd:101:8  */
  assign dp_readena = n6988_o; // (signal)
  /* ../../HW/src/top/cell.vhd:102:8  */
  assign dp_read_data_flow = n6989_o; // (signal)
  /* ../../HW/src/top/cell.vhd:103:8  */
  assign dp_read_stream = n6990_o; // (signal)
  /* ../../HW/src/top/cell.vhd:104:8  */
  assign dp_read_stream_id = n6991_o; // (signal)
  /* ../../HW/src/top/cell.vhd:105:8  */
  assign dp_read_data_type = n6992_o; // (signal)
  /* ../../HW/src/top/cell.vhd:106:8  */
  assign dp_read_gen_valid = n6993_o; // (signal)
  /* ../../HW/src/top/cell.vhd:107:8  */
  assign dp_readdata = n6996_o; // (signal)
  /* ../../HW/src/top/cell.vhd:108:8  */
  assign dp_readdata_vm = n6999_o; // (signal)
  /* ../../HW/src/top/cell.vhd:109:8  */
  assign dp_readena_r = n7000_q; // (signal)
  /* ../../HW/src/top/cell.vhd:110:8  */
  assign dp_readdata_r = n7001_q; // (signal)
  /* ../../HW/src/top/cell.vhd:111:8  */
  assign dp_readdata_vm_r = n7002_q; // (signal)
  /* ../../HW/src/top/cell.vhd:112:8  */
  assign dp_read_gen_valid_r = n7003_q; // (signal)
  /* ../../HW/src/top/cell.vhd:113:8  */
  assign dp_read_data_flow_r = n7004_q; // (signal)
  /* ../../HW/src/top/cell.vhd:114:8  */
  assign dp_read_data_type_r = n7005_q; // (signal)
  /* ../../HW/src/top/cell.vhd:115:8  */
  assign dp_read_stream_r = n7006_q; // (signal)
  /* ../../HW/src/top/cell.vhd:116:8  */
  assign dp_read_stream_id_r = n7007_q; // (signal)
  /* ../../HW/src/top/cell.vhd:117:8  */
  assign dp_read_vector = n7010_o; // (signal)
  /* ../../HW/src/top/cell.vhd:118:8  */
  assign dp_read_vector_r = n7011_q; // (signal)
  /* ../../HW/src/top/cell.vhd:119:8  */
  assign dp_read_vaddr = n7014_o; // (signal)
  /* ../../HW/src/top/cell.vhd:120:8  */
  assign dp_read_vaddr_r = n7015_q; // (signal)
  /* ../../HW/src/top/cell.vhd:122:8  */
  assign dp_rd_vm_in_r = n7016_q; // (signal)
  /* ../../HW/src/top/cell.vhd:123:8  */
  assign dp_wr_vm_in_r = n7017_q; // (signal)
  /* ../../HW/src/top/cell.vhd:124:8  */
  assign dp_code_in_r = n7018_q; // (signal)
  /* ../../HW/src/top/cell.vhd:125:8  */
  assign dp_rd_addr_in_r = n7019_q; // (signal)
  /* ../../HW/src/top/cell.vhd:126:8  */
  assign dp_rd_addr_step_in_r = n7020_q; // (signal)
  /* ../../HW/src/top/cell.vhd:127:8  */
  assign dp_rd_share_in_r = n7021_q; // (signal)
  /* ../../HW/src/top/cell.vhd:128:8  */
  assign dp_wr_addr_in_r = n7022_q; // (signal)
  /* ../../HW/src/top/cell.vhd:129:8  */
  assign dp_wr_addr_step_in_r = n7023_q; // (signal)
  /* ../../HW/src/top/cell.vhd:130:8  */
  assign dp_wr_fork_in_r = n7024_q; // (signal)
  /* ../../HW/src/top/cell.vhd:131:8  */
  assign dp_wr_share_in_r = n7025_q; // (signal)
  /* ../../HW/src/top/cell.vhd:132:8  */
  assign dp_wr_mcast_in_r = n7026_q; // (signal)
  /* ../../HW/src/top/cell.vhd:133:8  */
  assign dp_write_in_r = n7027_q; // (signal)
  /* ../../HW/src/top/cell.vhd:134:8  */
  assign dp_write_gen_valid_in_r = n7028_q; // (signal)
  /* ../../HW/src/top/cell.vhd:135:8  */
  assign dp_write_vector_in_r = n7029_q; // (signal)
  /* ../../HW/src/top/cell.vhd:136:8  */
  assign dp_write_scatter_in_r = n7030_q; // (signal)
  /* ../../HW/src/top/cell.vhd:137:8  */
  assign dp_read_in_r = n7031_q; // (signal)
  /* ../../HW/src/top/cell.vhd:138:8  */
  assign dp_rd_fork_in_r = n7032_q; // (signal)
  /* ../../HW/src/top/cell.vhd:139:8  */
  assign dp_read_vector_in_r = n7033_q; // (signal)
  /* ../../HW/src/top/cell.vhd:140:8  */
  assign dp_read_scatter_in_r = n7034_q; // (signal)
  /* ../../HW/src/top/cell.vhd:141:8  */
  assign dp_read_gen_valid_in_r = n7035_q; // (signal)
  /* ../../HW/src/top/cell.vhd:142:8  */
  assign dp_read_data_flow_in_r = n7036_q; // (signal)
  /* ../../HW/src/top/cell.vhd:143:8  */
  assign dp_read_data_type_in_r = n7037_q; // (signal)
  /* ../../HW/src/top/cell.vhd:144:8  */
  assign dp_read_stream_in_r = n7038_q; // (signal)
  /* ../../HW/src/top/cell.vhd:145:8  */
  assign dp_read_stream_id_in_r = n7039_q; // (signal)
  /* ../../HW/src/top/cell.vhd:146:8  */
  assign dp_writedata_in_r = n7040_q; // (signal)
  /* ../../HW/src/top/cell.vhd:147:8  */
  assign dp_config_in_r = n7041_q; // (signal)
  /* ../../HW/src/top/cell.vhd:170:16  */
  assign n6642_o = ~reset_in;
  /* ../../HW/src/top/cell.vhd:184:27  */
  assign n6645_o = dp_readena == 4'b0000;
  /* ../../HW/src/top/cell.vhd:184:13  */
  assign n6648_o = n6645_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/cell.vhd:189:48  */
  assign n6649_o = dp_readena & dp_read_gen_valid;
  /* ../../HW/src/top/cell.vhd:190:36  */
  assign n6651_o = n6649_o == 4'b0000;
  /* ../../HW/src/top/cell.vhd:190:13  */
  assign n6654_o = n6651_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n6655_o = dp_read_data_flow[1:0];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n6657_o = 2'b00 | n6655_o;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n6659_o = dp_read_data_flow[3:2];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n6660_o = n6657_o | n6659_o;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n6661_o = dp_read_data_flow[5:4];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n6662_o = n6660_o | n6661_o;
  /* ../../HW/src/top/cell.vhd:200:63  */
  assign n6663_o = dp_read_data_flow[7:6];
  /* ../../HW/src/top/cell.vhd:200:43  */
  assign n6664_o = n6662_o | n6663_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n6665_o = dp_read_stream[0];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n6667_o = 1'b0 | n6665_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n6669_o = dp_read_stream[1];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n6670_o = n6667_o | n6669_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n6671_o = dp_read_stream[2];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n6672_o = n6670_o | n6671_o;
  /* ../../HW/src/top/cell.vhd:206:54  */
  assign n6673_o = dp_read_stream[3];
  /* ../../HW/src/top/cell.vhd:206:37  */
  assign n6674_o = n6672_o | n6673_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n6675_o = dp_read_stream_id[1:0];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n6677_o = 2'b00 | n6675_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n6679_o = dp_read_stream_id[3:2];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n6680_o = n6677_o | n6679_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n6681_o = dp_read_stream_id[5:4];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n6682_o = n6680_o | n6681_o;
  /* ../../HW/src/top/cell.vhd:212:107  */
  assign n6683_o = dp_read_stream_id[7:6];
  /* ../../HW/src/top/cell.vhd:212:70  */
  assign n6684_o = n6682_o | n6683_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n6685_o = dp_read_data_type[1:0];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n6687_o = 2'b00 | n6685_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n6689_o = dp_read_data_type[3:2];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n6690_o = n6687_o | n6689_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n6691_o = dp_read_data_type[5:4];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n6692_o = n6690_o | n6691_o;
  /* ../../HW/src/top/cell.vhd:218:63  */
  assign n6693_o = dp_read_data_type[7:6];
  /* ../../HW/src/top/cell.vhd:218:43  */
  assign n6694_o = n6692_o | n6693_o;
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n6757_o = enable_in[0];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n1_gen1_pcore_i_n6758 = gen_reg_n1_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n1_gen1_pcore_i_n6759 = gen_reg_n1_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n1_gen1_pcore_i_n6760 = gen_reg_n1_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n1_gen1_pcore_i_n6761 = gen_reg_n1_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n1_gen1_pcore_i_n6762 = gen_reg_n1_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n1_gen1_pcore_i_n6763 = gen_reg_n1_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n1_gen1_pcore_i_n6764 = gen_reg_n1_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n1_gen1_pcore_i_n6765 = gen_reg_n1_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n1_gen1_pcore_i_n6766 = gen_reg_n1_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n1_gen1_pcore_i_n6767 = gen_reg_n1_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n1_gen1_pcore_i_n6768 = gen_reg_n1_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n1_gen1_pcore_i_n6769 = gen_reg_n1_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_0_0 gen_reg_n1_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n6757_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n1_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n1_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n1_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n1_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n1_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n1_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n1_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n1_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n1_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n1_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n1_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n1_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n6794_o = enable_in[1];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n2_gen1_pcore_i_n6795 = gen_reg_n2_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n2_gen1_pcore_i_n6796 = gen_reg_n2_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n2_gen1_pcore_i_n6797 = gen_reg_n2_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n2_gen1_pcore_i_n6798 = gen_reg_n2_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n2_gen1_pcore_i_n6799 = gen_reg_n2_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n2_gen1_pcore_i_n6800 = gen_reg_n2_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n2_gen1_pcore_i_n6801 = gen_reg_n2_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n2_gen1_pcore_i_n6802 = gen_reg_n2_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n2_gen1_pcore_i_n6803 = gen_reg_n2_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n2_gen1_pcore_i_n6804 = gen_reg_n2_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n2_gen1_pcore_i_n6805 = gen_reg_n2_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n2_gen1_pcore_i_n6806 = gen_reg_n2_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_0_1 gen_reg_n2_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n6794_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n2_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n2_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n2_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n2_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n2_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n2_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n2_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n2_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n2_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n2_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n2_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n2_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n6831_o = enable_in[2];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n3_gen1_pcore_i_n6832 = gen_reg_n3_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n3_gen1_pcore_i_n6833 = gen_reg_n3_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n3_gen1_pcore_i_n6834 = gen_reg_n3_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n3_gen1_pcore_i_n6835 = gen_reg_n3_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n3_gen1_pcore_i_n6836 = gen_reg_n3_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n3_gen1_pcore_i_n6837 = gen_reg_n3_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n3_gen1_pcore_i_n6838 = gen_reg_n3_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n3_gen1_pcore_i_n6839 = gen_reg_n3_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n3_gen1_pcore_i_n6840 = gen_reg_n3_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n3_gen1_pcore_i_n6841 = gen_reg_n3_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n3_gen1_pcore_i_n6842 = gen_reg_n3_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n3_gen1_pcore_i_n6843 = gen_reg_n3_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_0_2 gen_reg_n3_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n6831_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n3_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n3_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n3_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n3_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n3_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n3_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n3_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n3_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n3_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n3_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n3_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n3_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:254:31  */
  assign n6868_o = enable_in[3];
  /* ../../HW/src/top/cell.vhd:264:24  */
  assign gen_reg_n4_gen1_pcore_i_n6869 = gen_reg_n4_gen1_pcore_i_i_y_neg_out; // (signal)
  /* ../../HW/src/top/cell.vhd:265:25  */
  assign gen_reg_n4_gen1_pcore_i_n6870 = gen_reg_n4_gen1_pcore_i_i_y_zero_out; // (signal)
  /* ../../HW/src/top/cell.vhd:294:28  */
  assign gen_reg_n4_gen1_pcore_i_n6871 = gen_reg_n4_gen1_pcore_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/cell.vhd:295:31  */
  assign gen_reg_n4_gen1_pcore_i_n6872 = gen_reg_n4_gen1_pcore_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/cell.vhd:296:27  */
  assign gen_reg_n4_gen1_pcore_i_n6873 = gen_reg_n4_gen1_pcore_i_dp_readena_out; // (signal)
  /* ../../HW/src/top/cell.vhd:297:31  */
  assign gen_reg_n4_gen1_pcore_i_n6874 = gen_reg_n4_gen1_pcore_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/top/cell.vhd:298:30  */
  assign gen_reg_n4_gen1_pcore_i_n6875 = gen_reg_n4_gen1_pcore_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/top/cell.vhd:299:34  */
  assign gen_reg_n4_gen1_pcore_i_n6876 = gen_reg_n4_gen1_pcore_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/cell.vhd:300:33  */
  assign gen_reg_n4_gen1_pcore_i_n6877 = gen_reg_n4_gen1_pcore_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/top/cell.vhd:301:33  */
  assign gen_reg_n4_gen1_pcore_i_n6878 = gen_reg_n4_gen1_pcore_i_dp_read_data_type_out; // (signal)
  /* ../../HW/src/top/cell.vhd:302:31  */
  assign gen_reg_n4_gen1_pcore_i_n6879 = gen_reg_n4_gen1_pcore_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/top/cell.vhd:303:34  */
  assign gen_reg_n4_gen1_pcore_i_n6880 = gen_reg_n4_gen1_pcore_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/top/cell.vhd:236:1  */
  pcore_0_3 gen_reg_n4_gen1_pcore_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .instruction_mu_in(instruction_mu_in),
    .instruction_imu_in(instruction_imu_in),
    .instruction_mu_valid_in(instruction_mu_valid_in),
    .instruction_imu_valid_in(instruction_imu_valid_in),
    .vm_in(vm_in),
    .data_model_in(data_model_in),
    .enable_in(n6868_o),
    .tid_in(tid_in),
    .tid_valid1_in(tid_valid1_in),
    .pre_tid_in(pre_tid_in),
    .pre_tid_valid1_in(pre_tid_valid1_in),
    .pre_pre_tid_in(pre_pre_tid_in),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1_in),
    .pre_pre_vm_in(pre_pre_vm_in),
    .pre_pre_data_model_in(pre_pre_data_model_in),
    .pre_iregister_auto_in(pre_iregister_auto_in),
    .dp_rd_vm_in(dp_rd_vm_in_r),
    .dp_wr_vm_in(dp_wr_vm_in_r),
    .dp_code_in(dp_code_in_r),
    .dp_rd_addr_in(dp_rd_addr_in_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_in_r),
    .dp_rd_share_in(dp_rd_share_in_r),
    .dp_rd_fork_in(dp_rd_fork_in_r),
    .dp_wr_addr_in(dp_wr_addr_in_r),
    .dp_wr_addr_step_in(dp_wr_addr_step_in_r),
    .dp_wr_fork_in(dp_wr_fork_in_r),
    .dp_wr_share_in(dp_wr_share_in_r),
    .dp_wr_mcast_in(dp_wr_mcast_in_r),
    .dp_write_in(dp_write_in_r),
    .dp_write_gen_valid_in(dp_write_gen_valid_in_r),
    .dp_write_vector_in(dp_write_vector_in_r),
    .dp_write_scatter_in(dp_write_scatter_in_r),
    .dp_read_in(dp_read_in_r),
    .dp_read_vector_in(dp_read_vector_in_r),
    .dp_read_scatter_in(dp_read_scatter_in_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_in_r),
    .dp_read_data_flow_in(dp_read_data_flow_in_r),
    .dp_read_data_type_in(dp_read_data_type_in_r),
    .dp_read_stream_in(dp_read_stream_in_r),
    .dp_read_stream_id_in(dp_read_stream_id_in_r),
    .dp_writedata_in(dp_writedata_in_r),
    .dp_config_in_in(dp_config_in_r),
    .i_y_neg_out(gen_reg_n4_gen1_pcore_i_i_y_neg_out),
    .i_y_zero_out(gen_reg_n4_gen1_pcore_i_i_y_zero_out),
    .dp_readdata_out(gen_reg_n4_gen1_pcore_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_reg_n4_gen1_pcore_i_dp_readdata_vm_out),
    .dp_readena_out(gen_reg_n4_gen1_pcore_i_dp_readena_out),
    .dp_read_vector_out(gen_reg_n4_gen1_pcore_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_reg_n4_gen1_pcore_i_dp_read_vaddr_out),
    .dp_read_gen_valid_out(gen_reg_n4_gen1_pcore_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_reg_n4_gen1_pcore_i_dp_read_data_flow_out),
    .dp_read_data_type_out(gen_reg_n4_gen1_pcore_i_dp_read_data_type_out),
    .dp_read_stream_out(gen_reg_n4_gen1_pcore_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_reg_n4_gen1_pcore_i_dp_read_stream_id_out));
  /* ../../HW/src/top/cell.vhd:322:13  */
  assign n6907_o = ~reset_in;
  /* ../../HW/src/dp/dp.vhd:84:20  */
  assign n6988_o = {gen_reg_n4_gen1_pcore_i_n6873, gen_reg_n3_gen1_pcore_i_n6836, gen_reg_n2_gen1_pcore_i_n6799, gen_reg_n1_gen1_pcore_i_n6762};
  /* ../../HW/src/dp/dp.vhd:83:20  */
  assign n6989_o = {gen_reg_n4_gen1_pcore_i_n6877, gen_reg_n3_gen1_pcore_i_n6840, gen_reg_n2_gen1_pcore_i_n6803, gen_reg_n1_gen1_pcore_i_n6766};
  /* ../../HW/src/dp/dp.vhd:79:20  */
  assign n6990_o = {gen_reg_n4_gen1_pcore_i_n6879, gen_reg_n3_gen1_pcore_i_n6842, gen_reg_n2_gen1_pcore_i_n6805, gen_reg_n1_gen1_pcore_i_n6768};
  /* ../../HW/src/dp/dp.vhd:78:20  */
  assign n6991_o = {gen_reg_n4_gen1_pcore_i_n6880, gen_reg_n3_gen1_pcore_i_n6843, gen_reg_n2_gen1_pcore_i_n6806, gen_reg_n1_gen1_pcore_i_n6769};
  /* ../../HW/src/dp/dp.vhd:77:20  */
  assign n6992_o = {gen_reg_n4_gen1_pcore_i_n6878, gen_reg_n3_gen1_pcore_i_n6841, gen_reg_n2_gen1_pcore_i_n6804, gen_reg_n1_gen1_pcore_i_n6767};
  /* ../../HW/src/dp/dp.vhd:76:20  */
  assign n6993_o = {gen_reg_n4_gen1_pcore_i_n6876, gen_reg_n3_gen1_pcore_i_n6839, gen_reg_n2_gen1_pcore_i_n6802, gen_reg_n1_gen1_pcore_i_n6765};
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n6994_o = gen_reg_n1_gen1_pcore_i_n6760;
  assign n6994_o = gen_reg_n2_gen1_pcore_i_n6797;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n6995_o = n6994_o;
  assign n6995_o = gen_reg_n3_gen1_pcore_i_n6834;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n6996_o = n6995_o;
  assign n6996_o = gen_reg_n4_gen1_pcore_i_n6871;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n6997_o = gen_reg_n1_gen1_pcore_i_n6761;
  assign n6997_o = gen_reg_n2_gen1_pcore_i_n6798;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n6998_o = n6997_o;
  assign n6998_o = gen_reg_n3_gen1_pcore_i_n6835;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n6999_o = n6998_o;
  assign n6999_o = gen_reg_n4_gen1_pcore_i_n6872;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7000_q <= 1'b0;
    else
      n7000_q <= n6648_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7001_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n7001_q <= dp_readdata;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7002_q <= 1'b0;
    else
      n7002_q <= dp_readdata_vm;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7003_q <= 1'b0;
    else
      n7003_q <= n6654_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7004_q <= 2'b00;
    else
      n7004_q <= n6664_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7005_q <= 2'b00;
    else
      n7005_q <= n6694_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7006_q <= 1'b0;
    else
      n7006_q <= n6674_o;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7007_q <= 2'b00;
    else
      n7007_q <= n6684_o;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7008_o = gen_reg_n1_gen1_pcore_i_n6763;
  assign n7008_o = gen_reg_n2_gen1_pcore_i_n6800;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7009_o = n7008_o;
  assign n7009_o = gen_reg_n3_gen1_pcore_i_n6837;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7010_o = n7009_o;
  assign n7010_o = gen_reg_n4_gen1_pcore_i_n6874;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7011_q <= 3'b000;
    else
      n7011_q <= dp_read_vector;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7012_o = gen_reg_n1_gen1_pcore_i_n6764;
  assign n7012_o = gen_reg_n2_gen1_pcore_i_n6801;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7013_o = n7012_o;
  assign n7013_o = gen_reg_n3_gen1_pcore_i_n6838;
  /* ../../HW/src/top/cell.vhd:236:1  */
  assign n7014_o = n7013_o;
  assign n7014_o = gen_reg_n4_gen1_pcore_i_n6875;
  /* ../../HW/src/top/cell.vhd:182:9  */
  always @(posedge clock_in or posedge n6642_o)
    if (n6642_o)
      n7015_q <= 3'b000;
    else
      n7015_q <= dp_read_vaddr;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7016_q <= 1'b0;
    else
      n7016_q <= dp_rd_vm_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7017_q <= 1'b0;
    else
      n7017_q <= dp_wr_vm_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7018_q <= 1'b0;
    else
      n7018_q <= dp_code_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7019_q <= 22'b0000000000000000000000;
    else
      n7019_q <= dp_rd_addr_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7020_q <= 22'b0000000000000000000000;
    else
      n7020_q <= dp_rd_addr_step_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7021_q <= 1'b0;
    else
      n7021_q <= dp_rd_share_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7022_q <= 22'b0000000000000000000000;
    else
      n7022_q <= dp_wr_addr_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7023_q <= 22'b0000000000000000000000;
    else
      n7023_q <= dp_wr_addr_step_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7024_q <= 1'b0;
    else
      n7024_q <= dp_wr_fork_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7025_q <= 1'b0;
    else
      n7025_q <= dp_wr_share_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7026_q <= 6'b000000;
    else
      n7026_q <= dp_wr_mcast_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7027_q <= 1'b0;
    else
      n7027_q <= dp_write_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7028_q <= 1'b0;
    else
      n7028_q <= dp_write_gen_valid_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7029_q <= 3'b000;
    else
      n7029_q <= dp_write_vector_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7030_q <= 2'b00;
    else
      n7030_q <= dp_write_scatter_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7031_q <= 1'b0;
    else
      n7031_q <= dp_read_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7032_q <= 1'b0;
    else
      n7032_q <= dp_rd_fork_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7033_q <= 3'b000;
    else
      n7033_q <= dp_read_vector_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7034_q <= 2'b00;
    else
      n7034_q <= dp_read_scatter_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7035_q <= 1'b0;
    else
      n7035_q <= dp_read_gen_valid_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7036_q <= 2'b00;
    else
      n7036_q <= dp_read_data_flow_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7037_q <= 2'b00;
    else
      n7037_q <= dp_read_data_type_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7038_q <= 1'b0;
    else
      n7038_q <= dp_read_stream_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7039_q <= 2'b00;
    else
      n7039_q <= dp_read_stream_id_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7040_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n7040_q <= dp_writedata_in;
  /* ../../HW/src/top/cell.vhd:350:4  */
  always @(posedge clock_in or posedge n6907_o)
    if (n6907_o)
      n7041_q <= 1'b0;
    else
      n7041_q <= dp_config_in;
  /* ../../HW/src/top/cell.vhd:151:34  */
  assign n7042_o = dp_readena_r ? dp_readdata_r : 96'bz;
  /* ../../HW/src/top/cell.vhd:152:40  */
  assign n7043_o = dp_readena_r ? dp_readdata_vm_r : 1'bz;
  /* ../../HW/src/top/cell.vhd:159:40  */
  assign n7044_o = dp_readena_r ? dp_read_vector_r : 3'bz;
  /* ../../HW/src/top/cell.vhd:160:38  */
  assign n7045_o = dp_readena_r ? dp_read_vaddr_r : 3'bz;
  /* ../../HW/src/top/cell.vhd:154:46  */
  assign n7046_o = dp_readena_r ? dp_read_gen_valid_r : 1'bz;
  /* ../../HW/src/top/cell.vhd:155:46  */
  assign n7047_o = dp_readena_r ? dp_read_data_flow_r : 2'bz;
  /* ../../HW/src/top/cell.vhd:158:46  */
  assign n7048_o = dp_readena_r ? dp_read_data_type_r : 2'bz;
  /* ../../HW/src/top/cell.vhd:156:40  */
  assign n7049_o = dp_readena_r ? dp_read_stream_r : 1'bz;
  /* ../../HW/src/top/cell.vhd:157:46  */
  assign n7050_o = dp_readena_r ? dp_read_stream_id_r : 2'bz;
  /* ../../HW/src/top/cell.vhd:157:46  */
  assign n7051_o = {gen_reg_n4_gen1_pcore_i_n6869, gen_reg_n3_gen1_pcore_i_n6832, gen_reg_n2_gen1_pcore_i_n6795, gen_reg_n1_gen1_pcore_i_n6758};
  /* ../../HW/src/pcore/instr.vhd:216:5  */
  assign n7052_o = {gen_reg_n4_gen1_pcore_i_n6870, gen_reg_n3_gen1_pcore_i_n6833, gen_reg_n2_gen1_pcore_i_n6796, gen_reg_n1_gen1_pcore_i_n6759};
endmodule

module instr
  (input  clock_in,
   input  reset_in,
   input  dp_code_in,
   input  dp_config_in,
   input  [21:0] dp_wr_addr_in,
   input  dp_write_in,
   input  [95:0] dp_writedata_in,
   input  [7:0] i_y_neg_in,
   input  [7:0] i_y_zero_in,
   output [1:0] busy_out,
   output ready_out,
   output [79:0] instruction_mu_out,
   output [31:0] instruction_imu_out,
   output instruction_mu_valid_out,
   output instruction_imu_valid_out,
   output vm_out,
   output [1:0] data_model_out,
   output [7:0] enable_out,
   output [3:0] tid_out,
   output tid_valid1_out,
   output [3:0] pre_tid_out,
   output pre_tid_valid1_out,
   output [3:0] pre_pre_tid_out,
   output pre_pre_tid_valid1_out,
   output pre_pre_vm_out,
   output [1:0] pre_pre_data_model_out,
   output [27:0] pre_iregister_auto_out);
  wire [10:0] rom_addr;
  wire [10:0] rom_addr_plus_2;
  wire [127:0] rom_data;
  wire [63:0] instruction;
  wire instruction_write;
  wire instruction_write_r;
  wire [10:0] instruction_addr_r;
  wire [63:0] instruction_r;
  wire [10:0] task_start_addr_r;
  wire task_r;
  wire [4:0] task_pcore_max_r;
  wire task_vm_r;
  wire task_lockstep_r;
  wire [1:0] task_data_model_r;
  reg [3:0] task_tid_mask_r;
  wire [27:0] task_iregister_auto_r;
  wire y_neg_all;
  wire y_zero_all;
  wire dp_code_in_r;
  wire dp_config_in_r;
  wire [21:0] dp_wr_addr_in_r;
  wire dp_write_in_r;
  wire [95:0] dp_writedata_in_r;
  wire [63:0] n6359_o;
  wire n6361_o;
  wire n6362_o;
  wire n6366_o;
  wire n6367_o;
  wire n6371_o;
  wire n6372_o;
  wire [127:0] rom_i_n6374;
  wire [127:0] rom_i_instruction_out;
  wire [79:0] instr_fetch_i_n6377;
  wire [31:0] instr_fetch_i_n6378;
  wire instr_fetch_i_n6379;
  wire instr_fetch_i_n6380;
  wire instr_fetch_i_n6381;
  wire [1:0] instr_fetch_i_n6382;
  wire [3:0] instr_fetch_i_n6383;
  wire instr_fetch_i_n6384;
  wire [3:0] instr_fetch_i_n6385;
  wire instr_fetch_i_n6386;
  wire [3:0] instr_fetch_i_n6387;
  wire instr_fetch_i_n6388;
  wire instr_fetch_i_n6389;
  wire [1:0] instr_fetch_i_n6390;
  wire [7:0] instr_fetch_i_n6391;
  wire [27:0] instr_fetch_i_n6392;
  wire [10:0] instr_fetch_i_n6393;
  wire [10:0] instr_fetch_i_n6394;
  wire [1:0] instr_fetch_i_n6395;
  wire instr_fetch_i_n6396;
  wire [79:0] instr_fetch_i_instruction_mu_out;
  wire [31:0] instr_fetch_i_instruction_imu_out;
  wire instr_fetch_i_instruction_mu_valid_out;
  wire instr_fetch_i_instruction_imu_valid_out;
  wire instr_fetch_i_instruction_vm_out;
  wire [1:0] instr_fetch_i_instruction_data_model_out;
  wire [3:0] instr_fetch_i_instruction_tid_out;
  wire instr_fetch_i_instruction_tid_valid_out;
  wire [3:0] instr_fetch_i_instruction_pre_tid_out;
  wire instr_fetch_i_instruction_pre_tid_valid_out;
  wire [3:0] instr_fetch_i_instruction_pre_pre_tid_out;
  wire instr_fetch_i_instruction_pre_pre_tid_valid_out;
  wire instr_fetch_i_instruction_pre_pre_vm_out;
  wire [1:0] instr_fetch_i_instruction_pre_pre_data_model_out;
  wire [7:0] instr_fetch_i_instruction_pcore_enable_out;
  wire [27:0] instr_fetch_i_instruction_pre_iregister_auto_out;
  wire [10:0] instr_fetch_i_rom_addr_out;
  wire [10:0] instr_fetch_i_rom_addr_plus_2_out;
  wire [1:0] instr_fetch_i_busy_out;
  wire instr_fetch_i_ready_out;
  wire n6439_o;
  wire [10:0] n6441_o;
  wire n6462_o;
  wire [2:0] n6464_o;
  wire [10:0] n6465_o;
  wire [4:0] n6466_o;
  wire n6467_o;
  wire [3:0] n6468_o;
  wire [27:0] n6469_o;
  wire [1:0] n6470_o;
  wire n6472_o;
  wire n6475_o;
  wire n6476_o;
  wire n6478_o;
  wire n6480_o;
  wire n6481_o;
  wire n6482_o;
  wire n6485_o;
  wire [4:0] n6487_o;
  wire n6489_o;
  wire [1:0] n6491_o;
  wire [3:0] n6493_o;
  wire [27:0] n6495_o;
  reg n6572_q;
  reg [10:0] n6573_q;
  reg [63:0] n6574_q;
  reg [10:0] n6575_q;
  reg n6576_q;
  reg [4:0] n6577_q;
  reg n6578_q;
  reg n6579_q;
  reg [1:0] n6580_q;
  reg [3:0] n6581_q;
  reg [27:0] n6582_q;
  reg n6599_q;
  reg n6600_q;
  reg [21:0] n6601_q;
  reg n6602_q;
  reg [95:0] n6603_q;
  assign busy_out = instr_fetch_i_n6395;
  assign ready_out = instr_fetch_i_n6396;
  assign instruction_mu_out = instr_fetch_i_n6377;
  assign instruction_imu_out = instr_fetch_i_n6378;
  assign instruction_mu_valid_out = instr_fetch_i_n6379;
  assign instruction_imu_valid_out = instr_fetch_i_n6380;
  assign vm_out = instr_fetch_i_n6381;
  assign data_model_out = instr_fetch_i_n6382;
  assign enable_out = instr_fetch_i_n6391;
  assign tid_out = instr_fetch_i_n6383;
  assign tid_valid1_out = instr_fetch_i_n6384;
  assign pre_tid_out = instr_fetch_i_n6385;
  assign pre_tid_valid1_out = instr_fetch_i_n6386;
  assign pre_pre_tid_out = instr_fetch_i_n6387;
  assign pre_pre_tid_valid1_out = instr_fetch_i_n6388;
  assign pre_pre_vm_out = instr_fetch_i_n6389;
  assign pre_pre_data_model_out = instr_fetch_i_n6390;
  assign pre_iregister_auto_out = instr_fetch_i_n6392;
  /* ../../HW/src/pcore/instr.vhd:76:8  */
  assign rom_addr = instr_fetch_i_n6393; // (signal)
  /* ../../HW/src/pcore/instr.vhd:77:8  */
  assign rom_addr_plus_2 = instr_fetch_i_n6394; // (signal)
  /* ../../HW/src/pcore/instr.vhd:78:8  */
  assign rom_data = rom_i_n6374; // (signal)
  /* ../../HW/src/pcore/instr.vhd:80:8  */
  assign instruction = n6359_o; // (signal)
  /* ../../HW/src/pcore/instr.vhd:81:8  */
  assign instruction_write = n6362_o; // (signal)
  /* ../../HW/src/pcore/instr.vhd:82:8  */
  assign instruction_write_r = n6572_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:83:8  */
  assign instruction_addr_r = n6573_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:84:8  */
  assign instruction_r = n6574_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:88:8  */
  assign task_start_addr_r = n6575_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:89:8  */
  assign task_r = n6576_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:90:8  */
  assign task_pcore_max_r = n6577_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:91:8  */
  assign task_vm_r = n6578_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:92:8  */
  assign task_lockstep_r = n6579_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:93:8  */
  assign task_data_model_r = n6580_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:94:8  */
  always @*
    task_tid_mask_r = n6581_q; // (isignal)
  initial
    task_tid_mask_r = 4'b1111;
  /* ../../HW/src/pcore/instr.vhd:95:8  */
  assign task_iregister_auto_r = n6582_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:113:8  */
  assign y_neg_all = n6367_o; // (signal)
  /* ../../HW/src/pcore/instr.vhd:114:8  */
  assign y_zero_all = n6372_o; // (signal)
  /* ../../HW/src/pcore/instr.vhd:116:8  */
  assign dp_code_in_r = n6599_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:117:8  */
  assign dp_config_in_r = n6600_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:118:8  */
  assign dp_wr_addr_in_r = n6601_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:119:8  */
  assign dp_write_in_r = n6602_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:120:8  */
  assign dp_writedata_in_r = n6603_q; // (signal)
  /* ../../HW/src/pcore/instr.vhd:128:33  */
  assign n6359_o = dp_writedata_in_r[63:0];
  /* ../../HW/src/pcore/instr.vhd:130:50  */
  assign n6361_o = dp_code_in_r & dp_write_in_r;
  /* ../../HW/src/pcore/instr.vhd:130:26  */
  assign n6362_o = n6361_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr.vhd:132:33  */
  assign n6366_o = i_y_neg_in == 8'b00000000;
  /* ../../HW/src/pcore/instr.vhd:132:18  */
  assign n6367_o = n6366_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr.vhd:134:35  */
  assign n6371_o = i_y_zero_in == 8'b00000000;
  /* ../../HW/src/pcore/instr.vhd:134:19  */
  assign n6372_o = n6371_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr.vhd:140:38  */
  assign rom_i_n6374 = rom_i_instruction_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:136:1  */
  rom rom_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .rdaddress_in(rom_addr),
    .rdaddress_plus_2_in(rom_addr_plus_2),
    .wren_in(instruction_write_r),
    .wraddress_in(instruction_addr_r),
    .wrdata_in(instruction_r),
    .instruction_out(rom_i_instruction_out));
  /* ../../HW/src/pcore/instr.vhd:148:59  */
  assign instr_fetch_i_n6377 = instr_fetch_i_instruction_mu_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:149:60  */
  assign instr_fetch_i_n6378 = instr_fetch_i_instruction_imu_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:150:65  */
  assign instr_fetch_i_n6379 = instr_fetch_i_instruction_mu_valid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:151:66  */
  assign instr_fetch_i_n6380 = instr_fetch_i_instruction_imu_valid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:152:57  */
  assign instr_fetch_i_n6381 = instr_fetch_i_instruction_vm_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:153:117  */
  assign instr_fetch_i_n6382 = instr_fetch_i_instruction_data_model_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:154:59  */
  assign instr_fetch_i_n6383 = instr_fetch_i_instruction_tid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:155:65  */
  assign instr_fetch_i_n6384 = instr_fetch_i_instruction_tid_valid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:157:63  */
  assign instr_fetch_i_n6385 = instr_fetch_i_instruction_pre_tid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:158:69  */
  assign instr_fetch_i_n6386 = instr_fetch_i_instruction_pre_tid_valid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:159:67  */
  assign instr_fetch_i_n6387 = instr_fetch_i_instruction_pre_pre_tid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:160:73  */
  assign instr_fetch_i_n6388 = instr_fetch_i_instruction_pre_pre_tid_valid_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:162:67  */
  assign instr_fetch_i_n6389 = instr_fetch_i_instruction_pre_pre_vm_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:163:75  */
  assign instr_fetch_i_n6390 = instr_fetch_i_instruction_pre_pre_data_model_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:167:69  */
  assign instr_fetch_i_n6391 = instr_fetch_i_instruction_pcore_enable_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:165:75  */
  assign instr_fetch_i_n6392 = instr_fetch_i_instruction_pre_iregister_auto_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:172:51  */
  assign instr_fetch_i_n6393 = instr_fetch_i_rom_addr_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:173:58  */
  assign instr_fetch_i_n6394 = instr_fetch_i_rom_addr_plus_2_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:176:47  */
  assign instr_fetch_i_n6395 = instr_fetch_i_busy_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:177:48  */
  assign instr_fetch_i_n6396 = instr_fetch_i_ready_out; // (signal)
  /* ../../HW/src/pcore/instr.vhd:146:1  */
  instr_fetch instr_fetch_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .rom_data_in(rom_data),
    .task_start_addr_in(task_start_addr_r),
    .task_in(task_r),
    .task_pcore_max_in(task_pcore_max_r),
    .task_vm_in(task_vm_r),
    .task_lockstep_in(task_lockstep_r),
    .task_tid_mask_in(task_tid_mask_r),
    .task_iregister_auto_in(task_iregister_auto_r),
    .task_data_model_in(task_data_model_r),
    .i_y_neg_in(y_neg_all),
    .i_y_zero_in(y_zero_all),
    .instruction_mu_out(instr_fetch_i_instruction_mu_out),
    .instruction_imu_out(instr_fetch_i_instruction_imu_out),
    .instruction_mu_valid_out(instr_fetch_i_instruction_mu_valid_out),
    .instruction_imu_valid_out(instr_fetch_i_instruction_imu_valid_out),
    .instruction_vm_out(instr_fetch_i_instruction_vm_out),
    .instruction_data_model_out(instr_fetch_i_instruction_data_model_out),
    .instruction_tid_out(instr_fetch_i_instruction_tid_out),
    .instruction_tid_valid_out(instr_fetch_i_instruction_tid_valid_out),
    .instruction_pre_tid_out(instr_fetch_i_instruction_pre_tid_out),
    .instruction_pre_tid_valid_out(instr_fetch_i_instruction_pre_tid_valid_out),
    .instruction_pre_pre_tid_out(instr_fetch_i_instruction_pre_pre_tid_out),
    .instruction_pre_pre_tid_valid_out(instr_fetch_i_instruction_pre_pre_tid_valid_out),
    .instruction_pre_pre_vm_out(instr_fetch_i_instruction_pre_pre_vm_out),
    .instruction_pre_pre_data_model_out(instr_fetch_i_instruction_pre_pre_data_model_out),
    .instruction_pcore_enable_out(instr_fetch_i_instruction_pcore_enable_out),
    .instruction_pre_iregister_auto_out(instr_fetch_i_instruction_pre_iregister_auto_out),
    .rom_addr_out(instr_fetch_i_rom_addr_out),
    .rom_addr_plus_2_out(instr_fetch_i_rom_addr_plus_2_out),
    .busy_out(instr_fetch_i_busy_out),
    .ready_out(instr_fetch_i_ready_out));
  /* ../../HW/src/pcore/instr.vhd:189:16  */
  assign n6439_o = ~reset_in;
  /* ../../HW/src/pcore/instr.vhd:196:49  */
  assign n6441_o = dp_wr_addr_in_r[10:0];
  /* ../../HW/src/pcore/instr.vhd:216:16  */
  assign n6462_o = ~reset_in;
  /* ../../HW/src/pcore/instr.vhd:239:55  */
  assign n6464_o = dp_wr_addr_in_r[2:0];
  /* ../../HW/src/pcore/instr.vhd:241:50  */
  assign n6465_o = dp_writedata_in_r[10:0];
  /* ../../HW/src/pcore/instr.vhd:243:54  */
  assign n6466_o = dp_writedata_in_r[15:11];
  /* ../../HW/src/pcore/instr.vhd:245:43  */
  assign n6467_o = dp_writedata_in_r[16];
  /* ../../HW/src/pcore/instr.vhd:247:43  */
  assign n6468_o = dp_writedata_in_r[20:17];
  /* ../../HW/src/pcore/instr.vhd:249:58  */
  assign n6469_o = dp_writedata_in_r[48:21];
  /* ../../HW/src/pcore/instr.vhd:251:45  */
  assign n6470_o = dp_writedata_in_r[50:49];
  /* ../../HW/src/pcore/instr.vhd:253:30  */
  assign n6472_o = n6464_o == 3'b000;
  /* ../../HW/src/pcore/instr.vhd:253:12  */
  assign n6475_o = n6472_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/instr.vhd:258:34  */
  assign n6476_o = dp_config_in_r & dp_write_in_r;
  /* ../../HW/src/pcore/instr.vhd:258:78  */
  assign n6478_o = n6464_o == 3'b000;
  /* ../../HW/src/pcore/instr.vhd:258:123  */
  assign n6480_o = n6464_o == 3'b001;
  /* ../../HW/src/pcore/instr.vhd:258:104  */
  assign n6481_o = n6478_o | n6480_o;
  /* ../../HW/src/pcore/instr.vhd:258:57  */
  assign n6482_o = n6481_o & n6476_o;
  /* ../../HW/src/pcore/instr.vhd:258:12  */
  assign n6485_o = n6482_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/instr.vhd:258:12  */
  assign n6487_o = n6482_o ? n6466_o : 5'b00000;
  /* ../../HW/src/pcore/instr.vhd:258:12  */
  assign n6489_o = n6482_o ? n6467_o : 1'b0;
  /* ../../HW/src/pcore/instr.vhd:258:12  */
  assign n6491_o = n6482_o ? n6470_o : 2'b00;
  /* ../../HW/src/pcore/instr.vhd:258:12  */
  assign n6493_o = n6482_o ? n6468_o : 4'b1111;
  /* ../../HW/src/pcore/instr.vhd:258:12  */
  assign n6495_o = n6482_o ? n6469_o : 28'b0000000000000000000000000000;
  /* ../../HW/src/pcore/instr.vhd:194:9  */
  always @(posedge clock_in or posedge n6439_o)
    if (n6439_o)
      n6572_q <= 1'b0;
    else
      n6572_q <= instruction_write;
  /* ../../HW/src/pcore/instr.vhd:194:9  */
  always @(posedge clock_in or posedge n6439_o)
    if (n6439_o)
      n6573_q <= 11'b00000000000;
    else
      n6573_q <= n6441_o;
  /* ../../HW/src/pcore/instr.vhd:194:9  */
  always @(posedge clock_in or posedge n6439_o)
    if (n6439_o)
      n6574_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n6574_q <= instruction;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6575_q <= 11'b00000000000;
    else
      n6575_q <= n6465_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6576_q <= 1'b0;
    else
      n6576_q <= n6485_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6577_q <= 5'b00000;
    else
      n6577_q <= n6487_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6578_q <= 1'b0;
    else
      n6578_q <= n6475_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6579_q <= 1'b0;
    else
      n6579_q <= n6489_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6580_q <= 2'b00;
    else
      n6580_q <= n6491_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6581_q <= 4'b1111;
    else
      n6581_q <= n6493_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6582_q <= 28'b0000000000000000000000000000;
    else
      n6582_q <= n6495_o;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6599_q <= 1'b0;
    else
      n6599_q <= dp_code_in;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6600_q <= 1'b0;
    else
      n6600_q <= dp_config_in;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6601_q <= 22'b0000000000000000000000;
    else
      n6601_q <= dp_wr_addr_in;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6602_q <= 1'b0;
    else
      n6602_q <= dp_write_in;
  /* ../../HW/src/pcore/instr.vhd:231:9  */
  always @(posedge clock_in or posedge n6462_o)
    if (n6462_o)
      n6603_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n6603_q <= dp_writedata_in;
endmodule

module stream
  (input  clock_in,
   input  reset_in,
   input  [1:0] stream_id_in,
   input  [11:0] input_in,
   input  config_in,
   input  [8:0] config_reg_in,
   input  [23:0] config_data_in,
   output [11:0] output_out);
  wire [8:0] waddr_r;
  wire [8:0] \input ;
  wire [8:0] address;
  wire [23:0] writedata;
  wire [23:0] writedata_r;
  wire [23:0] y_mul;
  wire [23:0] y_mul_r;
  wire wena_r;
  wire [11:0] readdata2_r;
  wire [23:0] readdata_lookup;
  wire [23:0] readdata;
  wire [11:0] readdata_r;
  wire [11:0] readdata_rr;
  wire [4:0] remainder;
  wire [11:0] remainder_r;
  wire [11:0] remainder_rr;
  wire [11:0] \output ;
  wire [11:0] output_r;
  wire [12:0] y_mul_inc;
  wire [11:0] y_mul_round;
  wire [23:0] lookup_i_n6247;
  wire [23:0] lookup_i_q_a;
  wire [23:0] mul_i_n6250;
  wire [23:0] mul_i_z_out;
  wire [12:0] n6253_o;
  wire [12:0] n6255_o;
  wire [11:0] n6256_o;
  localparam n6257_o = 1'b1;
  wire [11:0] adder_i_n6258;
  wire [11:0] adder_i_z_out;
  wire [6:0] n6261_o;
  wire [8:0] n6262_o;
  wire [8:0] n6263_o;
  wire [4:0] n6264_o;
  wire n6270_o;
  wire [11:0] n6273_o;
  wire [11:0] n6274_o;
  wire n6279_o;
  wire [11:0] n6290_o;
  wire [8:0] n6326_o;
  reg [8:0] n6327_q;
  wire [23:0] n6328_o;
  reg [23:0] n6329_q;
  reg [23:0] n6330_q;
  reg n6331_q;
  reg [11:0] n6332_q;
  reg [11:0] n6333_q;
  reg [11:0] n6334_q;
  reg [11:0] n6336_q;
  reg [11:0] n6337_q;
  reg [11:0] n6339_q;
  assign output_out = output_r;
  /* ../../HW/src/pcore/stream.vhd:78:8  */
  assign waddr_r = n6327_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:79:8  */
  assign \input  = n6262_o; // (signal)
  /* ../../HW/src/pcore/stream.vhd:80:8  */
  assign address = n6263_o; // (signal)
  /* ../../HW/src/pcore/stream.vhd:81:8  */
  assign writedata = writedata_r; // (signal)
  /* ../../HW/src/pcore/stream.vhd:82:8  */
  assign writedata_r = n6329_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:83:8  */
  assign y_mul = mul_i_n6250; // (signal)
  /* ../../HW/src/pcore/stream.vhd:84:8  */
  assign y_mul_r = n6330_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:85:8  */
  assign wena_r = n6331_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:86:8  */
  assign readdata2_r = n6332_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:87:8  */
  assign readdata_lookup = lookup_i_n6247; // (signal)
  /* ../../HW/src/pcore/stream.vhd:88:8  */
  assign readdata = readdata_lookup; // (signal)
  /* ../../HW/src/pcore/stream.vhd:89:8  */
  assign readdata_r = n6333_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:90:8  */
  assign readdata_rr = n6334_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:92:8  */
  assign remainder = n6264_o; // (signal)
  /* ../../HW/src/pcore/stream.vhd:93:8  */
  assign remainder_r = n6336_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:94:8  */
  assign remainder_rr = n6337_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:96:8  */
  assign \output  = adder_i_n6258; // (signal)
  /* ../../HW/src/pcore/stream.vhd:97:8  */
  assign output_r = n6339_q; // (signal)
  /* ../../HW/src/pcore/stream.vhd:98:8  */
  assign y_mul_inc = n6255_o; // (signal)
  /* ../../HW/src/pcore/stream.vhd:99:8  */
  assign y_mul_round = n6256_o; // (signal)
  /* ../../HW/src/pcore/stream.vhd:113:13  */
  assign lookup_i_n6247 = lookup_i_q_a; // (signal)
  /* ../../HW/src/pcore/stream.vhd:102:1  */
  spram_512_9_24 lookup_i (
    .address_a(address),
    .clock0(clock_in),
    .data_a(writedata),
    .wren_a(wena_r),
    .q_a(lookup_i_q_a));
  /* ../../HW/src/pcore/stream.vhd:128:16  */
  assign mul_i_n6250 = mul_i_z_out; // (signal)
  /* ../../HW/src/pcore/stream.vhd:116:1  */
  multiplier_12_5ba93c9db0cff93f52b521d7420e43f6eda2784f mul_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .x_in(readdata2_r),
    .y_in(remainder_rr),
    .z_out(mul_i_z_out));
  /* ../../HW/src/pcore/stream.vhd:131:30  */
  assign n6253_o = y_mul_r[16:4];
  /* ../../HW/src/pcore/stream.vhd:131:140  */
  assign n6255_o = n6253_o + 13'b0000000000001;
  /* ../../HW/src/pcore/stream.vhd:134:42  */
  assign n6256_o = y_mul_inc[12:1];
  /* ../../HW/src/pcore/stream.vhd:146:14  */
  assign adder_i_n6258 = adder_i_z_out; // (signal)
  /* ../../HW/src/pcore/stream.vhd:136:1  */
  adder_12 adder_i (
    .x_in(y_mul_round),
    .y_in(readdata_rr),
    .add_sub_in(n6257_o),
    .z_out(adder_i_z_out));
  /* ../../HW/src/pcore/stream.vhd:151:51  */
  assign n6261_o = input_in[11:5];
  /* ../../HW/src/pcore/stream.vhd:151:41  */
  assign n6262_o = {stream_id_in, n6261_o};
  /* ../../HW/src/pcore/stream.vhd:153:20  */
  assign n6263_o = wena_r ? waddr_r : \input ;
  /* ../../HW/src/pcore/stream.vhd:155:22  */
  assign n6264_o = input_in[4:0];
  /* ../../HW/src/pcore/stream.vhd:171:17  */
  assign n6270_o = ~reset_in;
  /* ../../HW/src/pcore/stream.vhd:196:36  */
  assign n6273_o = readdata[11:0];
  /* ../../HW/src/pcore/stream.vhd:197:35  */
  assign n6274_o = readdata[23:12];
  /* ../../HW/src/pcore/stream.vhd:200:13  */
  assign n6279_o = config_in ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp.vhd:1071:32  */
  assign n6290_o = {7'b0000000, remainder};
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  assign n6326_o = config_in ? config_reg_in : waddr_r;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6327_q <= 9'b000000000;
    else
      n6327_q <= n6326_o;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  assign n6328_o = config_in ? config_data_in : writedata_r;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6329_q <= 24'b000000000000000000000000;
    else
      n6329_q <= n6328_o;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6330_q <= 24'b000000000000000000000000;
    else
      n6330_q <= y_mul;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6331_q <= 1'b0;
    else
      n6331_q <= n6279_o;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6332_q <= 12'b000000000000;
    else
      n6332_q <= n6273_o;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6333_q <= 12'b000000000000;
    else
      n6333_q <= n6274_o;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6334_q <= 12'b000000000000;
    else
      n6334_q <= readdata_r;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6336_q <= 12'b000000000000;
    else
      n6336_q <= n6290_o;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6337_q <= 12'b000000000000;
    else
      n6337_q <= remainder_r;
  /* ../../HW/src/pcore/stream.vhd:187:9  */
  always @(posedge clock_in or posedge n6270_o)
    if (n6270_o)
      n6339_q <= 12'b000000000000;
    else
      n6339_q <= \output ;
endmodule

module dp_0_611cf22eded7b64824a5f5c8e04751a6c8c2392b
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [11:0] bus_waddr_in,
   input  [11:0] bus_raddr_in,
   input  bus_write_in,
   input  bus_read_in,
   input  [31:0] bus_writedata_in,
   input  readmaster1_readdatavalid_in,
   input  readmaster1_readdatavalid_vm_in,
   input  [63:0] readmaster1_readdata_in,
   input  readmaster1_wait_request_in,
   input  writemaster1_wait_request_in,
   input  [47:0] writemaster1_counter_in,
   input  readmaster2_readdatavalid_in,
   input  readmaster2_readdatavalid_vm_in,
   input  [63:0] readmaster2_readdata_in,
   input  readmaster2_wait_request_in,
   input  writemaster2_wait_request_in,
   input  [47:0] writemaster2_counter_in,
   input  readmaster3_readdatavalid_in,
   input  readmaster3_readdatavalid_vm_in,
   input  [63:0] readmaster3_readdata_in,
   input  readmaster3_wait_request_in,
   input  writemaster3_wait_request_in,
   input  [23:0] writemaster3_counter_in,
   input  [1:0] task_busy_in,
   input  task_ready_in,
   input  [71:0] bar_in,
   input  ddr_tx_busy_in,
   output [31:0] bus_readdata_out,
   output bus_readdatavalid_out,
   output bus_writewait_out,
   output bus_readwait_out,
   output [21:0] readmaster1_addr_out,
   output readmaster1_fork_out,
   output readmaster1_addr_mode_out,
   output readmaster1_cs_out,
   output readmaster1_read_out,
   output readmaster1_read_vm_out,
   output [1:0] readmaster1_read_data_flow_out,
   output readmaster1_read_stream_out,
   output [1:0] readmaster1_read_stream_id_out,
   output [2:0] readmaster1_read_vector_out,
   output [1:0] readmaster1_read_scatter_out,
   output [4:0] readmaster1_burstlen_out,
   output [1:0] readmaster1_bus_id_out,
   output [1:0] readmaster1_data_type_out,
   output [1:0] readmaster1_data_model_out,
   output [21:0] writemaster1_addr_out,
   output writemaster1_fork_out,
   output writemaster1_addr_mode_out,
   output writemaster1_vm_out,
   output [5:0] writemaster1_mcast_out,
   output writemaster1_cs_out,
   output writemaster1_write_out,
   output [1:0] writemaster1_write_data_flow_out,
   output [2:0] writemaster1_write_vector_out,
   output writemaster1_write_stream_out,
   output [1:0] writemaster1_write_stream_id_out,
   output [1:0] writemaster1_write_scatter_out,
   output [63:0] writemaster1_writedata_out,
   output [4:0] writemaster1_burstlen_out,
   output [1:0] writemaster1_bus_id_out,
   output [1:0] writemaster1_data_type_out,
   output [1:0] writemaster1_data_model_out,
   output writemaster1_thread_out,
   output [17:0] readmaster2_addr_out,
   output readmaster2_fork_out,
   output readmaster2_cs_out,
   output readmaster2_read_out,
   output readmaster2_read_vm_out,
   output [2:0] readmaster2_read_vector_out,
   output [1:0] readmaster2_read_scatter_out,
   output [4:0] readmaster2_burstlen_out,
   output [1:0] readmaster2_bus_id_out,
   output [17:0] writemaster2_addr_out,
   output writemaster2_vm_out,
   output writemaster2_fork_out,
   output writemaster2_cs_out,
   output writemaster2_write_out,
   output [2:0] writemaster2_write_vector_out,
   output [1:0] writemaster2_write_scatter_out,
   output [63:0] writemaster2_writedata_out,
   output [4:0] writemaster2_burstlen_out,
   output [1:0] writemaster2_bus_id_out,
   output writemaster2_thread_out,
   output [31:0] readmaster3_addr_out,
   output readmaster3_cs_out,
   output readmaster3_read_out,
   output readmaster3_read_vm_out,
   output [2:0] readmaster3_read_vector_out,
   output [1:0] readmaster3_read_scatter_out,
   output [3:0] readmaster3_read_start_out,
   output [3:0] readmaster3_read_end_out,
   output [4:0] readmaster3_burstlen_out,
   output [1:0] readmaster3_bus_id_out,
   output [15:0] readmaster3_filler_data_out,
   output [31:0] writemaster3_addr_out,
   output writemaster3_cs_out,
   output writemaster3_write_out,
   output writemaster3_vm_out,
   output [2:0] writemaster3_write_vector_out,
   output [1:0] writemaster3_write_scatter_out,
   output [3:0] writemaster3_write_end_out,
   output [63:0] writemaster3_writedata_out,
   output [4:0] writemaster3_burstlen_out,
   output [8:0] writemaster3_burstlen2_out,
   output [4:0] writemaster3_burstlen3_out,
   output [1:0] writemaster3_bus_id_out,
   output writemaster3_thread_out,
   output [10:0] task_start_addr_out,
   output task_out,
   output task_pending_out,
   output task_vm_out,
   output [4:0] task_pcore_out,
   output task_lockstep_out,
   output [3:0] task_tid_mask_out,
   output [27:0] task_iregister_auto_out,
   output [1:0] task_data_model_out,
   output indication_avail_out);
  wire [1:0] ready;
  wire [1:0] valid;
  wire [1619:0] instruction;
  wire [1619:0] pre_instruction;
  wire gen_pcore_src_valid;
  wire gen_pcore_vm;
  wire [31:0] gen_pcore_src_addr;
  wire gen_pcore_src_addr_mode;
  wire gen_pcore_src_eof;
  wire [4:0] gen_pcore_src_burstlen;
  wire [31:0] gen_pcore_dst_addr;
  wire gen_pcore_dst_addr_mode;
  wire [4:0] gen_pcore_dst_burstlen;
  wire [1:0] gen_pcore_bus_id_source;
  wire [1:0] gen_pcore_bus_id_dest;
  wire gen_pcore_busy_dest;
  wire [1:0] gen_pcore_data_type_source;
  wire [1:0] gen_pcore_data_type_dest;
  wire [1:0] gen_pcore_data_model_source;
  wire [1:0] gen_pcore_data_model_dest;
  wire gen_pcore_thread;
  wire [5:0] gen_pcore_mcast;
  wire gen_pcore_fork;
  wire [2:0] gen_pcore_src_vector;
  wire [2:0] gen_pcore_dst_vector;
  wire [1:0] gen_pcore_src_scatter;
  wire [1:0] gen_pcore_dst_scatter;
  wire [3:0] gen_pcore_src_start;
  wire [3:0] gen_pcore_src_end;
  wire [3:0] gen_pcore_dst_end;
  wire [63:0] gen_pcore_data;
  wire [1:0] gen_pcore_data_flow;
  wire gen_pcore_src_stream;
  wire gen_pcore_dest_stream;
  wire [1:0] gen_pcore_stream_id;
  wire gen_sram_src_valid;
  wire gen_sram_vm;
  wire [31:0] gen_sram_src_addr;
  wire gen_sram_src_addr_mode;
  wire gen_sram_src_eof;
  wire [4:0] gen_sram_src_burstlen;
  wire [31:0] gen_sram_dst_addr;
  wire gen_sram_dst_addr_mode;
  wire [4:0] gen_sram_dst_burstlen;
  wire [1:0] gen_sram_bus_id_source;
  wire [1:0] gen_sram_bus_id_dest;
  wire gen_sram_busy_dest;
  wire [1:0] gen_sram_data_type_source;
  wire [1:0] gen_sram_data_type_dest;
  wire [1:0] gen_sram_data_model_source;
  wire [1:0] gen_sram_data_model_dest;
  wire gen_sram_thread;
  wire [5:0] gen_sram_mcast;
  wire gen_sram_fork;
  wire [2:0] gen_sram_src_vector;
  wire [2:0] gen_sram_dst_vector;
  wire [1:0] gen_sram_src_scatter;
  wire [1:0] gen_sram_dst_scatter;
  wire [3:0] gen_sram_src_start;
  wire [3:0] gen_sram_src_end;
  wire [3:0] gen_sram_dst_end;
  wire [63:0] gen_sram_data;
  wire [1:0] gen_sram_data_flow;
  wire gen_sram_src_stream;
  wire gen_sram_dest_stream;
  wire [1:0] gen_sram_stream_id;
  wire gen_ddr_src_valid;
  wire gen_ddr_vm;
  wire [31:0] gen_ddr_src_addr;
  wire gen_ddr_src_addr_mode;
  wire gen_ddr_src_eof;
  wire [4:0] gen_ddr_src_burstlen;
  wire [31:0] gen_ddr_dst_addr;
  wire gen_ddr_dst_addr_mode;
  wire [4:0] gen_ddr_dst_burstlen;
  wire [1:0] gen_ddr_bus_id_source;
  wire [1:0] gen_ddr_bus_id_dest;
  wire gen_ddr_busy_dest;
  wire [1:0] gen_ddr_data_type_source;
  wire [1:0] gen_ddr_data_type_dest;
  wire [1:0] gen_ddr_data_model_source;
  wire [1:0] gen_ddr_data_model_dest;
  wire gen_ddr_thread;
  wire [5:0] gen_ddr_mcast;
  wire gen_ddr_fork;
  wire [2:0] gen_ddr_src_vector;
  wire [2:0] gen_ddr_dst_vector;
  wire [1:0] gen_ddr_src_scatter;
  wire [1:0] gen_ddr_dst_scatter;
  wire [3:0] gen_ddr_src_start;
  wire [3:0] gen_ddr_src_end;
  wire [3:0] gen_ddr_dst_end;
  wire [63:0] gen_ddr_data;
  wire [1:0] gen_ddr_data_flow;
  wire gen_ddr_src_stream;
  wire gen_ddr_dest_stream;
  wire [1:0] gen_ddr_stream_id;
  wire [2:0] wr_datavalid;
  wire [95:0] wr_addr;
  wire [2:0] wr_fork;
  wire [2:0] wr_addr_mode;
  wire [2:0] wr_src_vm;
  wire [191:0] wr_data;
  wire [191:0] wr_readdata;
  wire [2:0] wr_readdatavalid;
  wire [2:0] wr_readdatavalid_vm;
  wire [14:0] wr_burstlen;
  wire [5:0] wr_bus_id;
  wire [2:0] wr_thread;
  wire [5:0] wr_data_type;
  wire [5:0] wr_data_model;
  wire [17:0] wr_mcast;
  wire [2:0] waitreq;
  wire wr_full;
  wire [2:0] wr_req;
  wire [2:0] wr_req_p0_pending;
  wire [2:0] wr_req_p1_pending;
  wire wr_sram_full;
  wire [2:0] wr_sram_req;
  wire [2:0] wr_sram_req_p0_pending;
  wire [2:0] wr_sram_req_p1_pending;
  wire wr_ddr_full;
  wire [2:0] wr_ddr_req;
  wire [2:0] wr_ddr_req_p0_pending;
  wire [2:0] wr_ddr_req_p1_pending;
  wire indication_avail;
  wire [2:0] full;
  wire [14:0] wr_maxburstlen;
  wire [2:0] pcore_read_pending_p0;
  wire [2:0] sram_read_pending_p0;
  wire [2:0] ddr_read_pending_p0;
  wire [2:0] pcore_read_pending_p1;
  wire [2:0] sram_read_pending_p1;
  wire [2:0] ddr_read_pending_p1;
  wire [8:0] wr_vector;
  wire [8:0] wr_sram_vector;
  wire [8:0] wr_ddr_vector;
  wire [5:0] wr_scatter;
  wire [5:0] wr_sram_scatter;
  wire [5:0] wr_ddr_scatter;
  wire [11:0] wr_end;
  wire [11:0] wr_sram_end;
  wire [11:0] wr_ddr_end;
  wire [5:0] wr_data_flow;
  wire [5:0] wr_sram_data_flow;
  wire [5:0] wr_ddr_data_flow;
  wire [2:0] wr_stream;
  wire [5:0] wr_stream_id;
  wire [31:0] log1;
  wire log1_valid;
  wire [31:0] log2;
  wire log2_valid;
  wire [31:0] readmaster1_addr;
  wire [31:0] readmaster2_addr;
  wire [31:0] readmaster3_addr;
  wire [31:0] writemaster1_addr;
  wire [31:0] writemaster2_addr;
  wire [31:0] writemaster3_addr;
  wire [21:0] n5147_o;
  wire [17:0] n5148_o;
  wire [15:0] n5149_o;
  wire [21:0] n5150_o;
  wire [17:0] n5151_o;
  wire [31:0] dp_fetch_1_i_n5153;
  wire dp_fetch_1_i_n5154;
  wire dp_fetch_1_i_n5155;
  wire dp_fetch_1_i_n5156;
  wire [1:0] dp_fetch_1_i_n5157;
  wire [1619:0] dp_fetch_1_i_n5158;
  wire [1619:0] dp_fetch_1_i_n5159;
  wire [10:0] dp_fetch_1_i_n5160;
  wire dp_fetch_1_i_n5161;
  wire dp_fetch_1_i_n5162;
  wire dp_fetch_1_i_n5163;
  wire [4:0] dp_fetch_1_i_n5164;
  wire dp_fetch_1_i_n5165;
  wire [3:0] dp_fetch_1_i_n5166;
  wire [27:0] dp_fetch_1_i_n5167;
  wire [1:0] dp_fetch_1_i_n5168;
  wire dp_fetch_1_i_n5169;
  wire [31:0] dp_fetch_1_i_bus_readdata_out;
  wire dp_fetch_1_i_bus_readdatavalid_out;
  wire dp_fetch_1_i_bus_writewait_out;
  wire dp_fetch_1_i_bus_readwait_out;
  wire [1:0] dp_fetch_1_i_instruction_valid_out;
  wire [2:0] dp_fetch_1_i_instruction_out_opcode;
  wire [3:0] dp_fetch_1_i_instruction_out_condition;
  wire dp_fetch_1_i_instruction_out_vm;
  wire [775:0] dp_fetch_1_i_instruction_out_source;
  wire [1:0] dp_fetch_1_i_instruction_out_source_bus_id;
  wire [1:0] dp_fetch_1_i_instruction_out_source_data_type;
  wire [775:0] dp_fetch_1_i_instruction_out_dest;
  wire [1:0] dp_fetch_1_i_instruction_out_dest_bus_id;
  wire [1:0] dp_fetch_1_i_instruction_out_dest_data_type;
  wire [5:0] dp_fetch_1_i_instruction_out_mcast;
  wire [23:0] dp_fetch_1_i_instruction_out_count;
  wire [15:0] dp_fetch_1_i_instruction_out_data;
  wire dp_fetch_1_i_instruction_out_repeat;
  wire dp_fetch_1_i_instruction_out_source_addr_mode;
  wire dp_fetch_1_i_instruction_out_dest_addr_mode;
  wire dp_fetch_1_i_instruction_out_stream_process;
  wire [1:0] dp_fetch_1_i_instruction_out_stream_process_id;
  wire [2:0] dp_fetch_1_i_pre_instruction_out_opcode;
  wire [3:0] dp_fetch_1_i_pre_instruction_out_condition;
  wire dp_fetch_1_i_pre_instruction_out_vm;
  wire [775:0] dp_fetch_1_i_pre_instruction_out_source;
  wire [1:0] dp_fetch_1_i_pre_instruction_out_source_bus_id;
  wire [1:0] dp_fetch_1_i_pre_instruction_out_source_data_type;
  wire [775:0] dp_fetch_1_i_pre_instruction_out_dest;
  wire [1:0] dp_fetch_1_i_pre_instruction_out_dest_bus_id;
  wire [1:0] dp_fetch_1_i_pre_instruction_out_dest_data_type;
  wire [5:0] dp_fetch_1_i_pre_instruction_out_mcast;
  wire [23:0] dp_fetch_1_i_pre_instruction_out_count;
  wire [15:0] dp_fetch_1_i_pre_instruction_out_data;
  wire dp_fetch_1_i_pre_instruction_out_repeat;
  wire dp_fetch_1_i_pre_instruction_out_source_addr_mode;
  wire dp_fetch_1_i_pre_instruction_out_dest_addr_mode;
  wire dp_fetch_1_i_pre_instruction_out_stream_process;
  wire [1:0] dp_fetch_1_i_pre_instruction_out_stream_process_id;
  wire [10:0] dp_fetch_1_i_task_start_addr_out;
  wire dp_fetch_1_i_task_pending_out;
  wire dp_fetch_1_i_task_out;
  wire dp_fetch_1_i_task_vm_out;
  wire [4:0] dp_fetch_1_i_task_pcore_out;
  wire dp_fetch_1_i_task_lockstep_out;
  wire [3:0] dp_fetch_1_i_task_tid_mask_out;
  wire [27:0] dp_fetch_1_i_task_iregister_auto_out;
  wire [1:0] dp_fetch_1_i_task_data_model_out;
  wire dp_fetch_1_i_indication_avail_out;
  wire [1619:0] n5175_o;
  wire [1619:0] n5177_o;
  wire [1:0] dp_gen_core_i_n5206;
  wire [31:0] dp_gen_core_i_n5207;
  wire dp_gen_core_i_n5208;
  wire [31:0] dp_gen_core_i_n5209;
  wire dp_gen_core_i_n5210;
  wire dp_gen_core_i_n5211;
  wire dp_gen_core_i_n5212;
  wire dp_gen_core_i_n5213;
  wire [1:0] dp_gen_core_i_n5214;
  wire dp_gen_core_i_n5215;
  wire dp_gen_core_i_n5216;
  wire [1:0] dp_gen_core_i_n5217;
  wire [2:0] dp_gen_core_i_n5218;
  wire [2:0] dp_gen_core_i_n5219;
  wire [1:0] dp_gen_core_i_n5220;
  wire [1:0] dp_gen_core_i_n5221;
  wire [3:0] dp_gen_core_i_n5222;
  wire [3:0] dp_gen_core_i_n5223;
  wire [3:0] dp_gen_core_i_n5224;
  wire [31:0] dp_gen_core_i_n5225;
  wire dp_gen_core_i_n5226;
  wire [31:0] dp_gen_core_i_n5227;
  wire dp_gen_core_i_n5228;
  wire dp_gen_core_i_n5229;
  wire [1:0] dp_gen_core_i_n5230;
  wire [1:0] dp_gen_core_i_n5231;
  wire [1:0] dp_gen_core_i_n5232;
  wire [1:0] dp_gen_core_i_n5233;
  wire dp_gen_core_i_n5234;
  wire [1:0] dp_gen_core_i_n5235;
  wire [1:0] dp_gen_core_i_n5236;
  wire [4:0] dp_gen_core_i_n5237;
  wire [4:0] dp_gen_core_i_n5238;
  wire dp_gen_core_i_n5239;
  wire [5:0] dp_gen_core_i_n5240;
  wire [63:0] dp_gen_core_i_n5241;
  wire dp_gen_core_i_n5242;
  wire dp_gen_core_i_n5243;
  wire dp_gen_core_i_n5244;
  wire [1:0] dp_gen_core_i_n5245;
  wire dp_gen_core_i_n5246;
  wire dp_gen_core_i_n5247;
  wire [1:0] dp_gen_core_i_n5248;
  wire [2:0] dp_gen_core_i_n5249;
  wire [2:0] dp_gen_core_i_n5250;
  wire [1:0] dp_gen_core_i_n5251;
  wire [1:0] dp_gen_core_i_n5252;
  wire [3:0] dp_gen_core_i_n5253;
  wire [3:0] dp_gen_core_i_n5254;
  wire [3:0] dp_gen_core_i_n5255;
  wire [31:0] dp_gen_core_i_n5256;
  wire dp_gen_core_i_n5257;
  wire [31:0] dp_gen_core_i_n5258;
  wire dp_gen_core_i_n5259;
  wire dp_gen_core_i_n5260;
  wire [1:0] dp_gen_core_i_n5261;
  wire [1:0] dp_gen_core_i_n5262;
  wire [1:0] dp_gen_core_i_n5263;
  wire [1:0] dp_gen_core_i_n5264;
  wire dp_gen_core_i_n5265;
  wire [1:0] dp_gen_core_i_n5266;
  wire [1:0] dp_gen_core_i_n5267;
  wire [4:0] dp_gen_core_i_n5268;
  wire [4:0] dp_gen_core_i_n5269;
  wire dp_gen_core_i_n5270;
  wire [5:0] dp_gen_core_i_n5271;
  wire [63:0] dp_gen_core_i_n5272;
  wire dp_gen_core_i_n5273;
  wire dp_gen_core_i_n5274;
  wire dp_gen_core_i_n5275;
  wire [1:0] dp_gen_core_i_n5276;
  wire dp_gen_core_i_n5277;
  wire dp_gen_core_i_n5278;
  wire [1:0] dp_gen_core_i_n5279;
  wire [2:0] dp_gen_core_i_n5280;
  wire [2:0] dp_gen_core_i_n5281;
  wire [1:0] dp_gen_core_i_n5282;
  wire [1:0] dp_gen_core_i_n5283;
  wire [3:0] dp_gen_core_i_n5284;
  wire [3:0] dp_gen_core_i_n5285;
  wire [3:0] dp_gen_core_i_n5286;
  wire [31:0] dp_gen_core_i_n5287;
  wire dp_gen_core_i_n5288;
  wire [31:0] dp_gen_core_i_n5289;
  wire dp_gen_core_i_n5290;
  wire dp_gen_core_i_n5291;
  wire [1:0] dp_gen_core_i_n5292;
  wire [1:0] dp_gen_core_i_n5293;
  wire [1:0] dp_gen_core_i_n5294;
  wire [1:0] dp_gen_core_i_n5295;
  wire dp_gen_core_i_n5296;
  wire [1:0] dp_gen_core_i_n5297;
  wire [1:0] dp_gen_core_i_n5298;
  wire [4:0] dp_gen_core_i_n5299;
  wire [4:0] dp_gen_core_i_n5300;
  wire dp_gen_core_i_n5301;
  wire [5:0] dp_gen_core_i_n5302;
  wire [63:0] dp_gen_core_i_n5303;
  wire [1:0] dp_gen_core_i_ready_out;
  wire [31:0] dp_gen_core_i_log1_out;
  wire dp_gen_core_i_log1_valid_out;
  wire [31:0] dp_gen_core_i_log2_out;
  wire dp_gen_core_i_log2_valid_out;
  wire dp_gen_core_i_gen_pcore_src_valid_out;
  wire dp_gen_core_i_gen_pcore_vm_out;
  wire dp_gen_core_i_gen_pcore_fork_out;
  wire [1:0] dp_gen_core_i_gen_pcore_data_flow_out;
  wire dp_gen_core_i_gen_pcore_src_stream_out;
  wire dp_gen_core_i_gen_pcore_dest_stream_out;
  wire [1:0] dp_gen_core_i_gen_pcore_stream_id_out;
  wire [2:0] dp_gen_core_i_gen_pcore_src_vector_out;
  wire [2:0] dp_gen_core_i_gen_pcore_dst_vector_out;
  wire [1:0] dp_gen_core_i_gen_pcore_src_scatter_out;
  wire [1:0] dp_gen_core_i_gen_pcore_dst_scatter_out;
  wire [3:0] dp_gen_core_i_gen_pcore_src_start_out;
  wire [3:0] dp_gen_core_i_gen_pcore_src_end_out;
  wire [3:0] dp_gen_core_i_gen_pcore_dst_end_out;
  wire [31:0] dp_gen_core_i_gen_pcore_src_addr_out;
  wire dp_gen_core_i_gen_pcore_src_addr_mode_out;
  wire [31:0] dp_gen_core_i_gen_pcore_dst_addr_out;
  wire dp_gen_core_i_gen_pcore_dst_addr_mode_out;
  wire dp_gen_core_i_gen_pcore_src_eof_out;
  wire [1:0] dp_gen_core_i_gen_pcore_bus_id_source_out;
  wire [1:0] dp_gen_core_i_gen_pcore_data_type_source_out;
  wire [1:0] dp_gen_core_i_gen_pcore_data_model_source_out;
  wire [1:0] dp_gen_core_i_gen_pcore_bus_id_dest_out;
  wire dp_gen_core_i_gen_pcore_busy_dest_out;
  wire [1:0] dp_gen_core_i_gen_pcore_data_type_dest_out;
  wire [1:0] dp_gen_core_i_gen_pcore_data_model_dest_out;
  wire [4:0] dp_gen_core_i_gen_pcore_src_burstlen_out;
  wire [4:0] dp_gen_core_i_gen_pcore_dst_burstlen_out;
  wire dp_gen_core_i_gen_pcore_thread_out;
  wire [5:0] dp_gen_core_i_gen_pcore_mcast_out;
  wire [63:0] dp_gen_core_i_gen_pcore_data_out;
  wire dp_gen_core_i_gen_sram_src_valid_out;
  wire dp_gen_core_i_gen_sram_vm_out;
  wire dp_gen_core_i_gen_sram_fork_out;
  wire [1:0] dp_gen_core_i_gen_sram_data_flow_out;
  wire dp_gen_core_i_gen_sram_src_stream_out;
  wire dp_gen_core_i_gen_sram_dest_stream_out;
  wire [1:0] dp_gen_core_i_gen_sram_stream_id_out;
  wire [2:0] dp_gen_core_i_gen_sram_src_vector_out;
  wire [2:0] dp_gen_core_i_gen_sram_dst_vector_out;
  wire [1:0] dp_gen_core_i_gen_sram_src_scatter_out;
  wire [1:0] dp_gen_core_i_gen_sram_dst_scatter_out;
  wire [3:0] dp_gen_core_i_gen_sram_src_start_out;
  wire [3:0] dp_gen_core_i_gen_sram_src_end_out;
  wire [3:0] dp_gen_core_i_gen_sram_dst_end_out;
  wire [31:0] dp_gen_core_i_gen_sram_src_addr_out;
  wire dp_gen_core_i_gen_sram_src_addr_mode_out;
  wire [31:0] dp_gen_core_i_gen_sram_dst_addr_out;
  wire dp_gen_core_i_gen_sram_dst_addr_mode_out;
  wire dp_gen_core_i_gen_sram_src_eof_out;
  wire [1:0] dp_gen_core_i_gen_sram_bus_id_source_out;
  wire [1:0] dp_gen_core_i_gen_sram_data_type_source_out;
  wire [1:0] dp_gen_core_i_gen_sram_data_model_source_out;
  wire [1:0] dp_gen_core_i_gen_sram_bus_id_dest_out;
  wire dp_gen_core_i_gen_sram_busy_dest_out;
  wire [1:0] dp_gen_core_i_gen_sram_data_type_dest_out;
  wire [1:0] dp_gen_core_i_gen_sram_data_model_dest_out;
  wire [4:0] dp_gen_core_i_gen_sram_src_burstlen_out;
  wire [4:0] dp_gen_core_i_gen_sram_dst_burstlen_out;
  wire dp_gen_core_i_gen_sram_thread_out;
  wire [5:0] dp_gen_core_i_gen_sram_mcast_out;
  wire [63:0] dp_gen_core_i_gen_sram_data_out;
  wire dp_gen_core_i_gen_ddr_src_valid_out;
  wire dp_gen_core_i_gen_ddr_vm_out;
  wire dp_gen_core_i_gen_ddr_fork_out;
  wire [1:0] dp_gen_core_i_gen_ddr_data_flow_out;
  wire dp_gen_core_i_gen_ddr_src_stream_out;
  wire dp_gen_core_i_gen_ddr_dest_stream_out;
  wire [1:0] dp_gen_core_i_gen_ddr_stream_id_out;
  wire [2:0] dp_gen_core_i_gen_ddr_src_vector_out;
  wire [2:0] dp_gen_core_i_gen_ddr_dst_vector_out;
  wire [1:0] dp_gen_core_i_gen_ddr_src_scatter_out;
  wire [1:0] dp_gen_core_i_gen_ddr_dst_scatter_out;
  wire [3:0] dp_gen_core_i_gen_ddr_src_start_out;
  wire [3:0] dp_gen_core_i_gen_ddr_src_end_out;
  wire [3:0] dp_gen_core_i_gen_ddr_dst_end_out;
  wire [31:0] dp_gen_core_i_gen_ddr_src_addr_out;
  wire dp_gen_core_i_gen_ddr_src_addr_mode_out;
  wire [31:0] dp_gen_core_i_gen_ddr_dst_addr_out;
  wire dp_gen_core_i_gen_ddr_dst_addr_mode_out;
  wire dp_gen_core_i_gen_ddr_src_eof_out;
  wire [1:0] dp_gen_core_i_gen_ddr_bus_id_source_out;
  wire [1:0] dp_gen_core_i_gen_ddr_data_type_source_out;
  wire [1:0] dp_gen_core_i_gen_ddr_data_model_source_out;
  wire [1:0] dp_gen_core_i_gen_ddr_bus_id_dest_out;
  wire dp_gen_core_i_gen_ddr_busy_dest_out;
  wire [1:0] dp_gen_core_i_gen_ddr_data_type_dest_out;
  wire [1:0] dp_gen_core_i_gen_ddr_data_model_dest_out;
  wire [4:0] dp_gen_core_i_gen_ddr_src_burstlen_out;
  wire [4:0] dp_gen_core_i_gen_ddr_dst_burstlen_out;
  wire dp_gen_core_i_gen_ddr_thread_out;
  wire [5:0] dp_gen_core_i_gen_ddr_mcast_out;
  wire [63:0] dp_gen_core_i_gen_ddr_data_out;
  wire [2:0] n5305_o;
  wire [3:0] n5306_o;
  wire n5307_o;
  wire [775:0] n5308_o;
  wire [1:0] n5309_o;
  wire [1:0] n5310_o;
  wire [775:0] n5311_o;
  wire [1:0] n5312_o;
  wire [1:0] n5313_o;
  wire [5:0] n5314_o;
  wire [23:0] n5315_o;
  wire [15:0] n5316_o;
  wire n5317_o;
  wire n5318_o;
  wire n5319_o;
  wire n5320_o;
  wire [1:0] n5321_o;
  wire [2:0] n5322_o;
  wire [3:0] n5323_o;
  wire n5324_o;
  wire [775:0] n5325_o;
  wire [1:0] n5326_o;
  wire [1:0] n5327_o;
  wire [775:0] n5328_o;
  wire [1:0] n5329_o;
  wire [1:0] n5330_o;
  wire [5:0] n5331_o;
  wire [23:0] n5332_o;
  wire [15:0] n5333_o;
  wire n5334_o;
  wire n5335_o;
  wire n5336_o;
  wire n5337_o;
  wire [1:0] n5338_o;
  wire [31:0] dp_source1_i_n5534;
  wire dp_source1_i_n5535;
  wire dp_source1_i_n5536;
  wire dp_source1_i_n5537;
  wire dp_source1_i_n5538;
  wire dp_source1_i_n5539;
  wire [1:0] dp_source1_i_n5540;
  wire dp_source1_i_n5541;
  wire [1:0] dp_source1_i_n5542;
  wire [2:0] dp_source1_i_n5543;
  wire [1:0] dp_source1_i_n5544;
  wire [4:0] dp_source1_i_n5547;
  wire [1:0] dp_source1_i_n5548;
  wire [1:0] dp_source1_i_n5549;
  wire [1:0] dp_source1_i_n5550;
  wire dp_source1_i_n5551;
  wire [2:0] dp_source1_i_n5552;
  wire [2:0] dp_source1_i_n5553;
  wire [2:0] dp_source1_i_n5554;
  wire [2:0] n5555_o;
  wire [5:0] dp_source1_i_n5556;
  wire [8:0] dp_source1_i_n5557;
  wire [2:0] dp_source1_i_n5558;
  wire [5:0] dp_source1_i_n5559;
  wire [5:0] dp_source1_i_n5560;
  wire [11:0] dp_source1_i_n5561;
  wire [31:0] dp_source1_i_n5562;
  wire dp_source1_i_n5563;
  wire dp_source1_i_n5564;
  wire dp_source1_i_n5565;
  wire dp_source1_i_n5566;
  wire [63:0] dp_source1_i_n5567;
  wire dp_source1_i_n5568;
  wire dp_source1_i_n5569;
  wire [63:0] dp_source1_i_n5570;
  wire [4:0] dp_source1_i_n5571;
  wire [1:0] dp_source1_i_n5572;
  wire dp_source1_i_n5573;
  wire [1:0] dp_source1_i_n5574;
  wire [1:0] dp_source1_i_n5575;
  wire [5:0] dp_source1_i_n5576;
  wire [31:0] dp_source1_i_bus_addr_out;
  wire dp_source1_i_bus_addr_mode_out;
  wire dp_source1_i_bus_cs_out;
  wire dp_source1_i_bus_read_out;
  wire dp_source1_i_bus_read_vm_out;
  wire dp_source1_i_bus_read_fork_out;
  wire [1:0] dp_source1_i_bus_read_data_flow_out;
  wire dp_source1_i_bus_read_stream_out;
  wire [1:0] dp_source1_i_bus_read_stream_id_out;
  wire [2:0] dp_source1_i_bus_read_vector_out;
  wire [1:0] dp_source1_i_bus_read_scatter_out;
  wire [3:0] dp_source1_i_bus_read_start_out;
  wire [3:0] dp_source1_i_bus_read_end_out;
  wire [4:0] dp_source1_i_bus_burstlen_out;
  wire [1:0] dp_source1_i_bus_id_out;
  wire [1:0] dp_source1_i_bus_data_type_out;
  wire [1:0] dp_source1_i_bus_data_model_out;
  wire dp_source1_i_gen_waitreq_out;
  wire [2:0] dp_source1_i_wr_req_out;
  wire [2:0] dp_source1_i_wr_req_pending_p0_out;
  wire [2:0] dp_source1_i_wr_req_pending_p1_out;
  wire [5:0] dp_source1_i_wr_data_flow_out;
  wire [8:0] dp_source1_i_wr_vector_out;
  wire [2:0] dp_source1_i_wr_stream_out;
  wire [5:0] dp_source1_i_wr_stream_id_out;
  wire [5:0] dp_source1_i_wr_scatter_out;
  wire [11:0] dp_source1_i_wr_end_out;
  wire [31:0] dp_source1_i_wr_addr_out;
  wire dp_source1_i_wr_fork_out;
  wire dp_source1_i_wr_addr_mode_out;
  wire dp_source1_i_wr_src_vm_out;
  wire dp_source1_i_wr_datavalid_out;
  wire [63:0] dp_source1_i_wr_data_out;
  wire dp_source1_i_wr_readdatavalid_out;
  wire dp_source1_i_wr_readdatavalid_vm_out;
  wire [63:0] dp_source1_i_wr_readdata_out;
  wire [4:0] dp_source1_i_wr_burstlen_out;
  wire [1:0] dp_source1_i_wr_bus_id_out;
  wire dp_source1_i_wr_thread_out;
  wire [1:0] dp_source1_i_wr_data_type_out;
  wire [1:0] dp_source1_i_wr_data_model_out;
  wire [5:0] dp_source1_i_wr_mcast_out;
  wire n5636_o;
  wire n5637_o;
  wire n5638_o;
  wire n5640_o;
  wire n5641_o;
  wire n5642_o;
  wire n5644_o;
  wire n5645_o;
  wire n5646_o;
  wire [1:0] n5648_o;
  wire [1:0] n5649_o;
  wire [1:0] n5650_o;
  wire [2:0] n5652_o;
  wire [2:0] n5653_o;
  wire [2:0] n5654_o;
  wire n5656_o;
  wire [1:0] n5660_o;
  wire [1:0] n5664_o;
  wire [1:0] n5665_o;
  wire [1:0] n5666_o;
  wire [3:0] n5668_o;
  wire [3:0] n5669_o;
  wire [3:0] n5670_o;
  wire [31:0] dp_source2_i_n5686;
  wire dp_source2_i_n5688;
  wire dp_source2_i_n5689;
  wire dp_source2_i_n5690;
  wire dp_source2_i_n5691;
  wire [2:0] dp_source2_i_n5695;
  wire [1:0] dp_source2_i_n5696;
  wire [4:0] dp_source2_i_n5699;
  wire [1:0] dp_source2_i_n5700;
  wire dp_source2_i_n5703;
  wire [2:0] dp_source2_i_n5704;
  wire [2:0] dp_source2_i_n5705;
  wire [2:0] dp_source2_i_n5706;
  wire [2:0] n5707_o;
  wire [5:0] dp_source2_i_n5708;
  wire [8:0] dp_source2_i_n5709;
  wire [2:0] dp_source2_i_n5710;
  wire [5:0] dp_source2_i_n5711;
  wire [5:0] dp_source2_i_n5712;
  wire [11:0] dp_source2_i_n5713;
  wire [31:0] dp_source2_i_n5714;
  wire dp_source2_i_n5715;
  wire dp_source2_i_n5716;
  wire dp_source2_i_n5717;
  wire dp_source2_i_n5718;
  wire [63:0] dp_source2_i_n5719;
  wire dp_source2_i_n5720;
  wire dp_source2_i_n5721;
  wire [63:0] dp_source2_i_n5722;
  wire [4:0] dp_source2_i_n5723;
  wire [1:0] dp_source2_i_n5724;
  wire dp_source2_i_n5725;
  wire [1:0] dp_source2_i_n5726;
  wire [1:0] dp_source2_i_n5727;
  wire [5:0] dp_source2_i_n5728;
  wire [31:0] dp_source2_i_bus_addr_out;
  wire dp_source2_i_bus_addr_mode_out;
  wire dp_source2_i_bus_cs_out;
  wire dp_source2_i_bus_read_out;
  wire dp_source2_i_bus_read_vm_out;
  wire dp_source2_i_bus_read_fork_out;
  wire [1:0] dp_source2_i_bus_read_data_flow_out;
  wire dp_source2_i_bus_read_stream_out;
  wire [1:0] dp_source2_i_bus_read_stream_id_out;
  wire [2:0] dp_source2_i_bus_read_vector_out;
  wire [1:0] dp_source2_i_bus_read_scatter_out;
  wire [3:0] dp_source2_i_bus_read_start_out;
  wire [3:0] dp_source2_i_bus_read_end_out;
  wire [4:0] dp_source2_i_bus_burstlen_out;
  wire [1:0] dp_source2_i_bus_id_out;
  wire [1:0] dp_source2_i_bus_data_type_out;
  wire [1:0] dp_source2_i_bus_data_model_out;
  wire dp_source2_i_gen_waitreq_out;
  wire [2:0] dp_source2_i_wr_req_out;
  wire [2:0] dp_source2_i_wr_req_pending_p0_out;
  wire [2:0] dp_source2_i_wr_req_pending_p1_out;
  wire [5:0] dp_source2_i_wr_data_flow_out;
  wire [8:0] dp_source2_i_wr_vector_out;
  wire [2:0] dp_source2_i_wr_stream_out;
  wire [5:0] dp_source2_i_wr_stream_id_out;
  wire [5:0] dp_source2_i_wr_scatter_out;
  wire [11:0] dp_source2_i_wr_end_out;
  wire [31:0] dp_source2_i_wr_addr_out;
  wire dp_source2_i_wr_fork_out;
  wire dp_source2_i_wr_addr_mode_out;
  wire dp_source2_i_wr_src_vm_out;
  wire dp_source2_i_wr_datavalid_out;
  wire [63:0] dp_source2_i_wr_data_out;
  wire dp_source2_i_wr_readdatavalid_out;
  wire dp_source2_i_wr_readdatavalid_vm_out;
  wire [63:0] dp_source2_i_wr_readdata_out;
  wire [4:0] dp_source2_i_wr_burstlen_out;
  wire [1:0] dp_source2_i_wr_bus_id_out;
  wire dp_source2_i_wr_thread_out;
  wire [1:0] dp_source2_i_wr_data_type_out;
  wire [1:0] dp_source2_i_wr_data_model_out;
  wire [5:0] dp_source2_i_wr_mcast_out;
  wire n5782_o;
  wire n5783_o;
  wire n5784_o;
  wire n5786_o;
  wire n5787_o;
  wire n5788_o;
  wire n5790_o;
  wire n5791_o;
  wire n5792_o;
  wire [1:0] n5794_o;
  wire [1:0] n5795_o;
  wire [1:0] n5796_o;
  wire [2:0] n5798_o;
  wire [2:0] n5799_o;
  wire [2:0] n5800_o;
  wire n5802_o;
  wire [1:0] n5806_o;
  wire [1:0] n5810_o;
  wire [1:0] n5811_o;
  wire [1:0] n5812_o;
  wire [3:0] n5814_o;
  wire [3:0] n5815_o;
  wire [3:0] n5816_o;
  wire [31:0] dp_source3_i0_n5832;
  wire dp_source3_i0_n5834;
  wire dp_source3_i0_n5835;
  wire dp_source3_i0_n5836;
  wire [2:0] dp_source3_i0_n5841;
  wire [1:0] dp_source3_i0_n5842;
  wire [3:0] dp_source3_i0_n5843;
  wire [3:0] dp_source3_i0_n5844;
  wire [4:0] dp_source3_i0_n5845;
  wire [1:0] dp_source3_i0_n5846;
  wire dp_source3_i0_n5849;
  wire [2:0] dp_source3_i0_n5850;
  wire [2:0] dp_source3_i0_n5851;
  wire [2:0] dp_source3_i0_n5852;
  wire [2:0] n5853_o;
  wire [5:0] dp_source3_i0_n5854;
  wire [8:0] dp_source3_i0_n5855;
  wire [2:0] dp_source3_i0_n5856;
  wire [5:0] dp_source3_i0_n5857;
  wire [5:0] dp_source3_i0_n5858;
  wire [11:0] dp_source3_i0_n5859;
  wire [31:0] dp_source3_i0_n5860;
  wire dp_source3_i0_n5861;
  wire dp_source3_i0_n5862;
  wire dp_source3_i0_n5863;
  wire dp_source3_i0_n5864;
  wire [63:0] dp_source3_i0_n5865;
  wire dp_source3_i0_n5866;
  wire dp_source3_i0_n5867;
  wire [63:0] dp_source3_i0_n5868;
  wire [4:0] dp_source3_i0_n5869;
  wire [1:0] dp_source3_i0_n5870;
  wire dp_source3_i0_n5871;
  wire [1:0] dp_source3_i0_n5872;
  wire [1:0] dp_source3_i0_n5873;
  wire [5:0] dp_source3_i0_n5874;
  wire [31:0] dp_source3_i0_bus_addr_out;
  wire dp_source3_i0_bus_addr_mode_out;
  wire dp_source3_i0_bus_cs_out;
  wire dp_source3_i0_bus_read_out;
  wire dp_source3_i0_bus_read_vm_out;
  wire dp_source3_i0_bus_read_fork_out;
  wire [1:0] dp_source3_i0_bus_read_data_flow_out;
  wire dp_source3_i0_bus_read_stream_out;
  wire [1:0] dp_source3_i0_bus_read_stream_id_out;
  wire [2:0] dp_source3_i0_bus_read_vector_out;
  wire [1:0] dp_source3_i0_bus_read_scatter_out;
  wire [3:0] dp_source3_i0_bus_read_start_out;
  wire [3:0] dp_source3_i0_bus_read_end_out;
  wire [4:0] dp_source3_i0_bus_burstlen_out;
  wire [1:0] dp_source3_i0_bus_id_out;
  wire [1:0] dp_source3_i0_bus_data_type_out;
  wire [1:0] dp_source3_i0_bus_data_model_out;
  wire dp_source3_i0_gen_waitreq_out;
  wire [2:0] dp_source3_i0_wr_req_out;
  wire [2:0] dp_source3_i0_wr_req_pending_p0_out;
  wire [2:0] dp_source3_i0_wr_req_pending_p1_out;
  wire [5:0] dp_source3_i0_wr_data_flow_out;
  wire [8:0] dp_source3_i0_wr_vector_out;
  wire [2:0] dp_source3_i0_wr_stream_out;
  wire [5:0] dp_source3_i0_wr_stream_id_out;
  wire [5:0] dp_source3_i0_wr_scatter_out;
  wire [11:0] dp_source3_i0_wr_end_out;
  wire [31:0] dp_source3_i0_wr_addr_out;
  wire dp_source3_i0_wr_fork_out;
  wire dp_source3_i0_wr_addr_mode_out;
  wire dp_source3_i0_wr_src_vm_out;
  wire dp_source3_i0_wr_datavalid_out;
  wire [63:0] dp_source3_i0_wr_data_out;
  wire dp_source3_i0_wr_readdatavalid_out;
  wire dp_source3_i0_wr_readdatavalid_vm_out;
  wire [63:0] dp_source3_i0_wr_readdata_out;
  wire [4:0] dp_source3_i0_wr_burstlen_out;
  wire [1:0] dp_source3_i0_wr_bus_id_out;
  wire dp_source3_i0_wr_thread_out;
  wire [1:0] dp_source3_i0_wr_data_type_out;
  wire [1:0] dp_source3_i0_wr_data_model_out;
  wire [5:0] dp_source3_i0_wr_mcast_out;
  wire n5929_o;
  wire n5930_o;
  wire n5931_o;
  wire n5933_o;
  wire n5934_o;
  wire n5935_o;
  wire n5937_o;
  wire n5938_o;
  wire n5939_o;
  wire [1:0] n5941_o;
  wire [1:0] n5942_o;
  wire [1:0] n5943_o;
  wire [2:0] n5945_o;
  wire [2:0] n5946_o;
  wire [2:0] n5947_o;
  wire n5949_o;
  wire [1:0] n5953_o;
  wire [1:0] n5957_o;
  wire [1:0] n5958_o;
  wire [1:0] n5959_o;
  wire [3:0] n5961_o;
  wire [3:0] n5962_o;
  wire [3:0] n5963_o;
  wire [31:0] dp_sink1_i_n5979;
  wire dp_sink1_i_n5980;
  wire dp_sink1_i_n5981;
  wire dp_sink1_i_n5982;
  wire [1:0] dp_sink1_i_n5983;
  wire [2:0] dp_sink1_i_n5984;
  wire dp_sink1_i_n5985;
  wire [1:0] dp_sink1_i_n5986;
  wire [1:0] dp_sink1_i_n5987;
  wire [5:0] dp_sink1_i_n5989;
  wire dp_sink1_i_n5990;
  wire dp_sink1_i_n5991;
  wire [63:0] dp_sink1_i_n5992;
  wire [4:0] dp_sink1_i_n5993;
  wire [1:0] dp_sink1_i_n5996;
  wire [1:0] dp_sink1_i_n5997;
  wire [1:0] dp_sink1_i_n5998;
  wire dp_sink1_i_n5999;
  wire [4:0] dp_sink1_i_n6000;
  wire dp_sink1_i_n6001;
  wire [2:0] dp_sink1_i_n6002;
  wire [2:0] dp_sink1_i_n6003;
  wire [31:0] dp_sink1_i_bus_addr_out;
  wire dp_sink1_i_bus_fork_out;
  wire dp_sink1_i_bus_addr_mode_out;
  wire dp_sink1_i_bus_vm_out;
  wire [1:0] dp_sink1_i_bus_data_flow_out;
  wire [2:0] dp_sink1_i_bus_vector_out;
  wire dp_sink1_i_bus_stream_out;
  wire [1:0] dp_sink1_i_bus_stream_id_out;
  wire [1:0] dp_sink1_i_bus_scatter_out;
  wire [3:0] dp_sink1_i_bus_end_out;
  wire [5:0] dp_sink1_i_bus_mcast_out;
  wire dp_sink1_i_bus_cs_out;
  wire dp_sink1_i_bus_write_out;
  wire [63:0] dp_sink1_i_bus_writedata_out;
  wire [4:0] dp_sink1_i_bus_burstlen_out;
  wire [8:0] dp_sink1_i_bus_burstlen2_out;
  wire [4:0] dp_sink1_i_bus_burstlen3_out;
  wire [1:0] dp_sink1_i_bus_id_out;
  wire [1:0] dp_sink1_i_bus_data_type_out;
  wire [1:0] dp_sink1_i_bus_data_model_out;
  wire dp_sink1_i_bus_thread_out;
  wire [4:0] dp_sink1_i_wr_maxburstlen_out;
  wire dp_sink1_i_wr_full_out;
  wire [2:0] dp_sink1_i_read_pending_p0_out;
  wire [2:0] dp_sink1_i_read_pending_p1_out;
  wire [31:0] dp_sink2_i_n6051;
  wire dp_sink2_i_n6052;
  wire dp_sink2_i_n6054;
  wire [2:0] dp_sink2_i_n6056;
  wire [1:0] dp_sink2_i_n6059;
  wire dp_sink2_i_n6062;
  wire dp_sink2_i_n6063;
  wire [63:0] dp_sink2_i_n6064;
  wire [4:0] dp_sink2_i_n6065;
  wire [1:0] dp_sink2_i_n6068;
  wire dp_sink2_i_n6071;
  wire [4:0] dp_sink2_i_n6072;
  wire dp_sink2_i_n6073;
  localparam [2:0] n6074_o = 3'b000;
  localparam [5:0] n6075_o = 6'b000000;
  wire [2:0] dp_sink2_i_n6076;
  wire [2:0] dp_sink2_i_n6077;
  wire [31:0] dp_sink2_i_bus_addr_out;
  wire dp_sink2_i_bus_fork_out;
  wire dp_sink2_i_bus_addr_mode_out;
  wire dp_sink2_i_bus_vm_out;
  wire [1:0] dp_sink2_i_bus_data_flow_out;
  wire [2:0] dp_sink2_i_bus_vector_out;
  wire dp_sink2_i_bus_stream_out;
  wire [1:0] dp_sink2_i_bus_stream_id_out;
  wire [1:0] dp_sink2_i_bus_scatter_out;
  wire [3:0] dp_sink2_i_bus_end_out;
  wire [5:0] dp_sink2_i_bus_mcast_out;
  wire dp_sink2_i_bus_cs_out;
  wire dp_sink2_i_bus_write_out;
  wire [63:0] dp_sink2_i_bus_writedata_out;
  wire [4:0] dp_sink2_i_bus_burstlen_out;
  wire [8:0] dp_sink2_i_bus_burstlen2_out;
  wire [4:0] dp_sink2_i_bus_burstlen3_out;
  wire [1:0] dp_sink2_i_bus_id_out;
  wire [1:0] dp_sink2_i_bus_data_type_out;
  wire [1:0] dp_sink2_i_bus_data_model_out;
  wire dp_sink2_i_bus_thread_out;
  wire [4:0] dp_sink2_i_wr_maxburstlen_out;
  wire dp_sink2_i_wr_full_out;
  wire [2:0] dp_sink2_i_read_pending_p0_out;
  wire [2:0] dp_sink2_i_read_pending_p1_out;
  wire [31:0] dp_sink3_i_n6118;
  wire dp_sink3_i_n6121;
  wire [2:0] dp_sink3_i_n6123;
  wire [1:0] dp_sink3_i_n6126;
  wire [3:0] dp_sink3_i_n6127;
  wire dp_sink3_i_n6129;
  wire dp_sink3_i_n6130;
  wire [63:0] dp_sink3_i_n6131;
  wire [4:0] dp_sink3_i_n6132;
  wire [8:0] dp_sink3_i_n6133;
  wire [4:0] dp_sink3_i_n6134;
  wire [1:0] dp_sink3_i_n6135;
  wire dp_sink3_i_n6138;
  wire [4:0] dp_sink3_i_n6139;
  wire dp_sink3_i_n6140;
  localparam [2:0] n6141_o = 3'b000;
  localparam [5:0] n6142_o = 6'b000000;
  wire [2:0] dp_sink3_i_n6143;
  wire [2:0] dp_sink3_i_n6144;
  wire [31:0] dp_sink3_i_bus_addr_out;
  wire dp_sink3_i_bus_fork_out;
  wire dp_sink3_i_bus_addr_mode_out;
  wire dp_sink3_i_bus_vm_out;
  wire [1:0] dp_sink3_i_bus_data_flow_out;
  wire [2:0] dp_sink3_i_bus_vector_out;
  wire dp_sink3_i_bus_stream_out;
  wire [1:0] dp_sink3_i_bus_stream_id_out;
  wire [1:0] dp_sink3_i_bus_scatter_out;
  wire [3:0] dp_sink3_i_bus_end_out;
  wire [5:0] dp_sink3_i_bus_mcast_out;
  wire dp_sink3_i_bus_cs_out;
  wire dp_sink3_i_bus_write_out;
  wire [63:0] dp_sink3_i_bus_writedata_out;
  wire [4:0] dp_sink3_i_bus_burstlen_out;
  wire [8:0] dp_sink3_i_bus_burstlen2_out;
  wire [4:0] dp_sink3_i_bus_burstlen3_out;
  wire [1:0] dp_sink3_i_bus_id_out;
  wire [1:0] dp_sink3_i_bus_data_type_out;
  wire [1:0] dp_sink3_i_bus_data_model_out;
  wire dp_sink3_i_bus_thread_out;
  wire [4:0] dp_sink3_i_wr_maxburstlen_out;
  wire dp_sink3_i_wr_full_out;
  wire [2:0] dp_sink3_i_read_pending_p0_out;
  wire [2:0] dp_sink3_i_read_pending_p1_out;
  wire [2:0] n6187_o;
  wire [95:0] n6188_o;
  wire [2:0] n6189_o;
  wire [2:0] n6190_o;
  wire [2:0] n6191_o;
  wire [191:0] n6192_o;
  wire [191:0] n6193_o;
  wire [2:0] n6194_o;
  wire [2:0] n6195_o;
  wire [14:0] n6196_o;
  wire [5:0] n6197_o;
  wire [2:0] n6198_o;
  wire [5:0] n6199_o;
  wire [5:0] n6200_o;
  wire [17:0] n6201_o;
  wire [2:0] n6202_o;
  wire [2:0] n6203_o;
  wire [2:0] n6204_o;
  wire [2:0] n6205_o;
  wire [2:0] n6206_o;
  wire [2:0] n6207_o;
  wire [2:0] n6208_o;
  wire [2:0] n6209_o;
  wire [2:0] n6210_o;
  wire [2:0] n6211_o;
  wire [2:0] n6226_o;
  wire [14:0] n6227_o;
  wire [8:0] n6228_o;
  wire [8:0] n6229_o;
  wire [8:0] n6230_o;
  wire [5:0] n6231_o;
  wire [5:0] n6232_o;
  wire [5:0] n6233_o;
  wire [11:0] n6234_o;
  wire [11:0] n6235_o;
  wire [11:0] n6236_o;
  wire [5:0] n6237_o;
  wire [5:0] n6238_o;
  wire [5:0] n6239_o;
  wire [2:0] n6240_o;
  wire [5:0] n6243_o;
  assign bus_readdata_out = dp_fetch_1_i_n5153;
  assign bus_readdatavalid_out = dp_fetch_1_i_n5154;
  assign bus_writewait_out = dp_fetch_1_i_n5155;
  assign bus_readwait_out = dp_fetch_1_i_n5156;
  assign readmaster1_addr_out = n5147_o;
  assign readmaster1_fork_out = dp_source1_i_n5539;
  assign readmaster1_addr_mode_out = dp_source1_i_n5535;
  assign readmaster1_cs_out = dp_source1_i_n5536;
  assign readmaster1_read_out = dp_source1_i_n5537;
  assign readmaster1_read_vm_out = dp_source1_i_n5538;
  assign readmaster1_read_data_flow_out = dp_source1_i_n5540;
  assign readmaster1_read_stream_out = dp_source1_i_n5541;
  assign readmaster1_read_stream_id_out = dp_source1_i_n5542;
  assign readmaster1_read_vector_out = dp_source1_i_n5543;
  assign readmaster1_read_scatter_out = dp_source1_i_n5544;
  assign readmaster1_burstlen_out = dp_source1_i_n5547;
  assign readmaster1_bus_id_out = dp_source1_i_n5548;
  assign readmaster1_data_type_out = dp_source1_i_n5549;
  assign readmaster1_data_model_out = dp_source1_i_n5550;
  assign writemaster1_addr_out = n5150_o;
  assign writemaster1_fork_out = dp_sink1_i_n5980;
  assign writemaster1_addr_mode_out = dp_sink1_i_n5981;
  assign writemaster1_vm_out = dp_sink1_i_n5982;
  assign writemaster1_mcast_out = dp_sink1_i_n5989;
  assign writemaster1_cs_out = dp_sink1_i_n5990;
  assign writemaster1_write_out = dp_sink1_i_n5991;
  assign writemaster1_write_data_flow_out = dp_sink1_i_n5983;
  assign writemaster1_write_vector_out = dp_sink1_i_n5984;
  assign writemaster1_write_stream_out = dp_sink1_i_n5985;
  assign writemaster1_write_stream_id_out = dp_sink1_i_n5986;
  assign writemaster1_write_scatter_out = dp_sink1_i_n5987;
  assign writemaster1_writedata_out = dp_sink1_i_n5992;
  assign writemaster1_burstlen_out = dp_sink1_i_n5993;
  assign writemaster1_bus_id_out = dp_sink1_i_n5996;
  assign writemaster1_data_type_out = dp_sink1_i_n5997;
  assign writemaster1_data_model_out = dp_sink1_i_n5998;
  assign writemaster1_thread_out = dp_sink1_i_n5999;
  assign readmaster2_addr_out = n5148_o;
  assign readmaster2_fork_out = dp_source2_i_n5691;
  assign readmaster2_cs_out = dp_source2_i_n5688;
  assign readmaster2_read_out = dp_source2_i_n5689;
  assign readmaster2_read_vm_out = dp_source2_i_n5690;
  assign readmaster2_read_vector_out = dp_source2_i_n5695;
  assign readmaster2_read_scatter_out = dp_source2_i_n5696;
  assign readmaster2_burstlen_out = dp_source2_i_n5699;
  assign readmaster2_bus_id_out = dp_source2_i_n5700;
  assign writemaster2_addr_out = n5151_o;
  assign writemaster2_vm_out = dp_sink2_i_n6054;
  assign writemaster2_fork_out = dp_sink2_i_n6052;
  assign writemaster2_cs_out = dp_sink2_i_n6062;
  assign writemaster2_write_out = dp_sink2_i_n6063;
  assign writemaster2_write_vector_out = dp_sink2_i_n6056;
  assign writemaster2_write_scatter_out = dp_sink2_i_n6059;
  assign writemaster2_writedata_out = dp_sink2_i_n6064;
  assign writemaster2_burstlen_out = dp_sink2_i_n6065;
  assign writemaster2_bus_id_out = dp_sink2_i_n6068;
  assign writemaster2_thread_out = dp_sink2_i_n6071;
  assign readmaster3_addr_out = readmaster3_addr;
  assign readmaster3_cs_out = dp_source3_i0_n5834;
  assign readmaster3_read_out = dp_source3_i0_n5835;
  assign readmaster3_read_vm_out = dp_source3_i0_n5836;
  assign readmaster3_read_vector_out = dp_source3_i0_n5841;
  assign readmaster3_read_scatter_out = dp_source3_i0_n5842;
  assign readmaster3_read_start_out = dp_source3_i0_n5843;
  assign readmaster3_read_end_out = dp_source3_i0_n5844;
  assign readmaster3_burstlen_out = dp_source3_i0_n5845;
  assign readmaster3_bus_id_out = dp_source3_i0_n5846;
  assign readmaster3_filler_data_out = n5149_o;
  assign writemaster3_addr_out = writemaster3_addr;
  assign writemaster3_cs_out = dp_sink3_i_n6129;
  assign writemaster3_write_out = dp_sink3_i_n6130;
  assign writemaster3_vm_out = dp_sink3_i_n6121;
  assign writemaster3_write_vector_out = dp_sink3_i_n6123;
  assign writemaster3_write_scatter_out = dp_sink3_i_n6126;
  assign writemaster3_write_end_out = dp_sink3_i_n6127;
  assign writemaster3_writedata_out = dp_sink3_i_n6131;
  assign writemaster3_burstlen_out = dp_sink3_i_n6132;
  assign writemaster3_burstlen2_out = dp_sink3_i_n6133;
  assign writemaster3_burstlen3_out = dp_sink3_i_n6134;
  assign writemaster3_bus_id_out = dp_sink3_i_n6135;
  assign writemaster3_thread_out = dp_sink3_i_n6138;
  assign task_start_addr_out = dp_fetch_1_i_n5160;
  assign task_out = dp_fetch_1_i_n5162;
  assign task_pending_out = dp_fetch_1_i_n5161;
  assign task_vm_out = dp_fetch_1_i_n5163;
  assign task_pcore_out = dp_fetch_1_i_n5164;
  assign task_lockstep_out = dp_fetch_1_i_n5165;
  assign task_tid_mask_out = dp_fetch_1_i_n5166;
  assign task_iregister_auto_out = dp_fetch_1_i_n5167;
  assign task_data_model_out = dp_fetch_1_i_n5168;
  assign indication_avail_out = indication_avail;
  /* ../../HW/src/dp/dp.vhd:200:8  */
  assign ready = dp_gen_core_i_n5206; // (signal)
  /* ../../HW/src/dp/dp.vhd:201:8  */
  assign valid = dp_fetch_1_i_n5157; // (signal)
  /* ../../HW/src/dp/dp.vhd:202:8  */
  assign instruction = dp_fetch_1_i_n5158; // (signal)
  /* ../../HW/src/dp/dp.vhd:203:8  */
  assign pre_instruction = dp_fetch_1_i_n5159; // (signal)
  /* ../../HW/src/dp/dp.vhd:205:8  */
  assign gen_pcore_src_valid = dp_gen_core_i_n5211; // (signal)
  /* ../../HW/src/dp/dp.vhd:206:8  */
  assign gen_pcore_vm = dp_gen_core_i_n5212; // (signal)
  /* ../../HW/src/dp/dp.vhd:207:8  */
  assign gen_pcore_src_addr = dp_gen_core_i_n5225; // (signal)
  /* ../../HW/src/dp/dp.vhd:208:8  */
  assign gen_pcore_src_addr_mode = dp_gen_core_i_n5226; // (signal)
  /* ../../HW/src/dp/dp.vhd:209:8  */
  assign gen_pcore_src_eof = dp_gen_core_i_n5229; // (signal)
  /* ../../HW/src/dp/dp.vhd:210:8  */
  assign gen_pcore_src_burstlen = dp_gen_core_i_n5237; // (signal)
  /* ../../HW/src/dp/dp.vhd:211:8  */
  assign gen_pcore_dst_addr = dp_gen_core_i_n5227; // (signal)
  /* ../../HW/src/dp/dp.vhd:212:8  */
  assign gen_pcore_dst_addr_mode = dp_gen_core_i_n5228; // (signal)
  /* ../../HW/src/dp/dp.vhd:213:8  */
  assign gen_pcore_dst_burstlen = dp_gen_core_i_n5238; // (signal)
  /* ../../HW/src/dp/dp.vhd:214:8  */
  assign gen_pcore_bus_id_source = dp_gen_core_i_n5230; // (signal)
  /* ../../HW/src/dp/dp.vhd:215:8  */
  assign gen_pcore_bus_id_dest = dp_gen_core_i_n5233; // (signal)
  /* ../../HW/src/dp/dp.vhd:216:8  */
  assign gen_pcore_busy_dest = dp_gen_core_i_n5234; // (signal)
  /* ../../HW/src/dp/dp.vhd:217:8  */
  assign gen_pcore_data_type_source = dp_gen_core_i_n5231; // (signal)
  /* ../../HW/src/dp/dp.vhd:218:8  */
  assign gen_pcore_data_type_dest = dp_gen_core_i_n5235; // (signal)
  /* ../../HW/src/dp/dp.vhd:219:8  */
  assign gen_pcore_data_model_source = dp_gen_core_i_n5232; // (signal)
  /* ../../HW/src/dp/dp.vhd:220:8  */
  assign gen_pcore_data_model_dest = dp_gen_core_i_n5236; // (signal)
  /* ../../HW/src/dp/dp.vhd:221:8  */
  assign gen_pcore_thread = dp_gen_core_i_n5239; // (signal)
  /* ../../HW/src/dp/dp.vhd:222:8  */
  assign gen_pcore_mcast = dp_gen_core_i_n5240; // (signal)
  /* ../../HW/src/dp/dp.vhd:223:8  */
  assign gen_pcore_fork = dp_gen_core_i_n5213; // (signal)
  /* ../../HW/src/dp/dp.vhd:224:8  */
  assign gen_pcore_src_vector = dp_gen_core_i_n5218; // (signal)
  /* ../../HW/src/dp/dp.vhd:225:8  */
  assign gen_pcore_dst_vector = dp_gen_core_i_n5219; // (signal)
  /* ../../HW/src/dp/dp.vhd:226:8  */
  assign gen_pcore_src_scatter = dp_gen_core_i_n5220; // (signal)
  /* ../../HW/src/dp/dp.vhd:227:8  */
  assign gen_pcore_dst_scatter = dp_gen_core_i_n5221; // (signal)
  /* ../../HW/src/dp/dp.vhd:228:8  */
  assign gen_pcore_src_start = dp_gen_core_i_n5222; // (signal)
  /* ../../HW/src/dp/dp.vhd:229:8  */
  assign gen_pcore_src_end = dp_gen_core_i_n5223; // (signal)
  /* ../../HW/src/dp/dp.vhd:230:8  */
  assign gen_pcore_dst_end = dp_gen_core_i_n5224; // (signal)
  /* ../../HW/src/dp/dp.vhd:231:8  */
  assign gen_pcore_data = dp_gen_core_i_n5241; // (signal)
  /* ../../HW/src/dp/dp.vhd:232:8  */
  assign gen_pcore_data_flow = dp_gen_core_i_n5214; // (signal)
  /* ../../HW/src/dp/dp.vhd:233:8  */
  assign gen_pcore_src_stream = dp_gen_core_i_n5215; // (signal)
  /* ../../HW/src/dp/dp.vhd:234:8  */
  assign gen_pcore_dest_stream = dp_gen_core_i_n5216; // (signal)
  /* ../../HW/src/dp/dp.vhd:235:8  */
  assign gen_pcore_stream_id = dp_gen_core_i_n5217; // (signal)
  /* ../../HW/src/dp/dp.vhd:237:8  */
  assign gen_sram_src_valid = dp_gen_core_i_n5242; // (signal)
  /* ../../HW/src/dp/dp.vhd:238:8  */
  assign gen_sram_vm = dp_gen_core_i_n5243; // (signal)
  /* ../../HW/src/dp/dp.vhd:239:8  */
  assign gen_sram_src_addr = dp_gen_core_i_n5256; // (signal)
  /* ../../HW/src/dp/dp.vhd:240:8  */
  assign gen_sram_src_addr_mode = dp_gen_core_i_n5257; // (signal)
  /* ../../HW/src/dp/dp.vhd:241:8  */
  assign gen_sram_src_eof = dp_gen_core_i_n5260; // (signal)
  /* ../../HW/src/dp/dp.vhd:242:8  */
  assign gen_sram_src_burstlen = dp_gen_core_i_n5268; // (signal)
  /* ../../HW/src/dp/dp.vhd:243:8  */
  assign gen_sram_dst_addr = dp_gen_core_i_n5258; // (signal)
  /* ../../HW/src/dp/dp.vhd:244:8  */
  assign gen_sram_dst_addr_mode = dp_gen_core_i_n5259; // (signal)
  /* ../../HW/src/dp/dp.vhd:245:8  */
  assign gen_sram_dst_burstlen = dp_gen_core_i_n5269; // (signal)
  /* ../../HW/src/dp/dp.vhd:246:8  */
  assign gen_sram_bus_id_source = dp_gen_core_i_n5261; // (signal)
  /* ../../HW/src/dp/dp.vhd:247:8  */
  assign gen_sram_bus_id_dest = dp_gen_core_i_n5264; // (signal)
  /* ../../HW/src/dp/dp.vhd:248:8  */
  assign gen_sram_busy_dest = dp_gen_core_i_n5265; // (signal)
  /* ../../HW/src/dp/dp.vhd:249:8  */
  assign gen_sram_data_type_source = dp_gen_core_i_n5262; // (signal)
  /* ../../HW/src/dp/dp.vhd:250:8  */
  assign gen_sram_data_type_dest = dp_gen_core_i_n5266; // (signal)
  /* ../../HW/src/dp/dp.vhd:251:8  */
  assign gen_sram_data_model_source = dp_gen_core_i_n5263; // (signal)
  /* ../../HW/src/dp/dp.vhd:252:8  */
  assign gen_sram_data_model_dest = dp_gen_core_i_n5267; // (signal)
  /* ../../HW/src/dp/dp.vhd:253:8  */
  assign gen_sram_thread = dp_gen_core_i_n5270; // (signal)
  /* ../../HW/src/dp/dp.vhd:254:8  */
  assign gen_sram_mcast = dp_gen_core_i_n5271; // (signal)
  /* ../../HW/src/dp/dp.vhd:255:8  */
  assign gen_sram_fork = dp_gen_core_i_n5244; // (signal)
  /* ../../HW/src/dp/dp.vhd:256:8  */
  assign gen_sram_src_vector = dp_gen_core_i_n5249; // (signal)
  /* ../../HW/src/dp/dp.vhd:257:8  */
  assign gen_sram_dst_vector = dp_gen_core_i_n5250; // (signal)
  /* ../../HW/src/dp/dp.vhd:258:8  */
  assign gen_sram_src_scatter = dp_gen_core_i_n5251; // (signal)
  /* ../../HW/src/dp/dp.vhd:259:8  */
  assign gen_sram_dst_scatter = dp_gen_core_i_n5252; // (signal)
  /* ../../HW/src/dp/dp.vhd:260:8  */
  assign gen_sram_src_start = dp_gen_core_i_n5253; // (signal)
  /* ../../HW/src/dp/dp.vhd:261:8  */
  assign gen_sram_src_end = dp_gen_core_i_n5254; // (signal)
  /* ../../HW/src/dp/dp.vhd:262:8  */
  assign gen_sram_dst_end = dp_gen_core_i_n5255; // (signal)
  /* ../../HW/src/dp/dp.vhd:263:8  */
  assign gen_sram_data = dp_gen_core_i_n5272; // (signal)
  /* ../../HW/src/dp/dp.vhd:264:8  */
  assign gen_sram_data_flow = dp_gen_core_i_n5245; // (signal)
  /* ../../HW/src/dp/dp.vhd:265:8  */
  assign gen_sram_src_stream = dp_gen_core_i_n5246; // (signal)
  /* ../../HW/src/dp/dp.vhd:266:8  */
  assign gen_sram_dest_stream = dp_gen_core_i_n5247; // (signal)
  /* ../../HW/src/dp/dp.vhd:267:8  */
  assign gen_sram_stream_id = dp_gen_core_i_n5248; // (signal)
  /* ../../HW/src/dp/dp.vhd:269:8  */
  assign gen_ddr_src_valid = dp_gen_core_i_n5273; // (signal)
  /* ../../HW/src/dp/dp.vhd:270:8  */
  assign gen_ddr_vm = dp_gen_core_i_n5274; // (signal)
  /* ../../HW/src/dp/dp.vhd:271:8  */
  assign gen_ddr_src_addr = dp_gen_core_i_n5287; // (signal)
  /* ../../HW/src/dp/dp.vhd:272:8  */
  assign gen_ddr_src_addr_mode = dp_gen_core_i_n5288; // (signal)
  /* ../../HW/src/dp/dp.vhd:273:8  */
  assign gen_ddr_src_eof = dp_gen_core_i_n5291; // (signal)
  /* ../../HW/src/dp/dp.vhd:274:8  */
  assign gen_ddr_src_burstlen = dp_gen_core_i_n5299; // (signal)
  /* ../../HW/src/dp/dp.vhd:275:8  */
  assign gen_ddr_dst_addr = dp_gen_core_i_n5289; // (signal)
  /* ../../HW/src/dp/dp.vhd:276:8  */
  assign gen_ddr_dst_addr_mode = dp_gen_core_i_n5290; // (signal)
  /* ../../HW/src/dp/dp.vhd:277:8  */
  assign gen_ddr_dst_burstlen = dp_gen_core_i_n5300; // (signal)
  /* ../../HW/src/dp/dp.vhd:278:8  */
  assign gen_ddr_bus_id_source = dp_gen_core_i_n5292; // (signal)
  /* ../../HW/src/dp/dp.vhd:279:8  */
  assign gen_ddr_bus_id_dest = dp_gen_core_i_n5295; // (signal)
  /* ../../HW/src/dp/dp.vhd:280:8  */
  assign gen_ddr_busy_dest = dp_gen_core_i_n5296; // (signal)
  /* ../../HW/src/dp/dp.vhd:281:8  */
  assign gen_ddr_data_type_source = dp_gen_core_i_n5293; // (signal)
  /* ../../HW/src/dp/dp.vhd:282:8  */
  assign gen_ddr_data_type_dest = dp_gen_core_i_n5297; // (signal)
  /* ../../HW/src/dp/dp.vhd:283:8  */
  assign gen_ddr_data_model_source = dp_gen_core_i_n5294; // (signal)
  /* ../../HW/src/dp/dp.vhd:284:8  */
  assign gen_ddr_data_model_dest = dp_gen_core_i_n5298; // (signal)
  /* ../../HW/src/dp/dp.vhd:285:8  */
  assign gen_ddr_thread = dp_gen_core_i_n5301; // (signal)
  /* ../../HW/src/dp/dp.vhd:286:8  */
  assign gen_ddr_mcast = dp_gen_core_i_n5302; // (signal)
  /* ../../HW/src/dp/dp.vhd:287:8  */
  assign gen_ddr_fork = dp_gen_core_i_n5275; // (signal)
  /* ../../HW/src/dp/dp.vhd:288:8  */
  assign gen_ddr_src_vector = dp_gen_core_i_n5280; // (signal)
  /* ../../HW/src/dp/dp.vhd:289:8  */
  assign gen_ddr_dst_vector = dp_gen_core_i_n5281; // (signal)
  /* ../../HW/src/dp/dp.vhd:290:8  */
  assign gen_ddr_src_scatter = dp_gen_core_i_n5282; // (signal)
  /* ../../HW/src/dp/dp.vhd:291:8  */
  assign gen_ddr_dst_scatter = dp_gen_core_i_n5283; // (signal)
  /* ../../HW/src/dp/dp.vhd:292:8  */
  assign gen_ddr_src_start = dp_gen_core_i_n5284; // (signal)
  /* ../../HW/src/dp/dp.vhd:293:8  */
  assign gen_ddr_src_end = dp_gen_core_i_n5285; // (signal)
  /* ../../HW/src/dp/dp.vhd:294:8  */
  assign gen_ddr_dst_end = dp_gen_core_i_n5286; // (signal)
  /* ../../HW/src/dp/dp.vhd:295:8  */
  assign gen_ddr_data = dp_gen_core_i_n5303; // (signal)
  /* ../../HW/src/dp/dp.vhd:296:8  */
  assign gen_ddr_data_flow = dp_gen_core_i_n5276; // (signal)
  /* ../../HW/src/dp/dp.vhd:297:8  */
  assign gen_ddr_src_stream = dp_gen_core_i_n5277; // (signal)
  /* ../../HW/src/dp/dp.vhd:298:8  */
  assign gen_ddr_dest_stream = dp_gen_core_i_n5278; // (signal)
  /* ../../HW/src/dp/dp.vhd:299:8  */
  assign gen_ddr_stream_id = dp_gen_core_i_n5279; // (signal)
  /* ../../HW/src/dp/dp.vhd:301:8  */
  assign wr_datavalid = n6187_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:302:8  */
  assign wr_addr = n6188_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:303:8  */
  assign wr_fork = n6189_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:304:8  */
  assign wr_addr_mode = n6190_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:305:8  */
  assign wr_src_vm = n6191_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:306:8  */
  assign wr_data = n6192_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:307:8  */
  assign wr_readdata = n6193_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:308:8  */
  assign wr_readdatavalid = n6194_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:309:8  */
  assign wr_readdatavalid_vm = n6195_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:310:8  */
  assign wr_burstlen = n6196_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:311:8  */
  assign wr_bus_id = n6197_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:312:8  */
  assign wr_thread = n6198_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:313:8  */
  assign wr_data_type = n6199_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:314:8  */
  assign wr_data_model = n6200_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:315:8  */
  assign wr_mcast = n6201_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:317:8  */
  assign waitreq = n6202_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:318:8  */
  assign wr_full = dp_sink1_i_n6001; // (signal)
  /* ../../HW/src/dp/dp.vhd:319:8  */
  assign wr_req = n6203_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:320:8  */
  assign wr_req_p0_pending = n6204_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:321:8  */
  assign wr_req_p1_pending = n6205_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:323:8  */
  assign wr_sram_full = dp_sink2_i_n6073; // (signal)
  /* ../../HW/src/dp/dp.vhd:324:8  */
  assign wr_sram_req = n6206_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:325:8  */
  assign wr_sram_req_p0_pending = n6207_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:326:8  */
  assign wr_sram_req_p1_pending = n6208_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:328:8  */
  assign wr_ddr_full = dp_sink3_i_n6140; // (signal)
  /* ../../HW/src/dp/dp.vhd:329:8  */
  assign wr_ddr_req = n6209_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:330:8  */
  assign wr_ddr_req_p0_pending = n6210_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:331:8  */
  assign wr_ddr_req_p1_pending = n6211_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:333:8  */
  assign indication_avail = dp_fetch_1_i_n5169; // (signal)
  /* ../../HW/src/dp/dp.vhd:353:8  */
  assign full = n6226_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:355:8  */
  assign wr_maxburstlen = n6227_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:357:8  */
  assign pcore_read_pending_p0 = dp_sink1_i_n6002; // (signal)
  /* ../../HW/src/dp/dp.vhd:358:8  */
  assign sram_read_pending_p0 = dp_sink2_i_n6076; // (signal)
  /* ../../HW/src/dp/dp.vhd:359:8  */
  assign ddr_read_pending_p0 = dp_sink3_i_n6143; // (signal)
  /* ../../HW/src/dp/dp.vhd:361:8  */
  assign pcore_read_pending_p1 = dp_sink1_i_n6003; // (signal)
  /* ../../HW/src/dp/dp.vhd:362:8  */
  assign sram_read_pending_p1 = dp_sink2_i_n6077; // (signal)
  /* ../../HW/src/dp/dp.vhd:363:8  */
  assign ddr_read_pending_p1 = dp_sink3_i_n6144; // (signal)
  /* ../../HW/src/dp/dp.vhd:366:8  */
  assign wr_vector = n6228_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:367:8  */
  assign wr_sram_vector = n6229_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:368:8  */
  assign wr_ddr_vector = n6230_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:369:8  */
  assign wr_scatter = n6231_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:370:8  */
  assign wr_sram_scatter = n6232_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:371:8  */
  assign wr_ddr_scatter = n6233_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:372:8  */
  assign wr_end = n6234_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:373:8  */
  assign wr_sram_end = n6235_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:374:8  */
  assign wr_ddr_end = n6236_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:376:8  */
  assign wr_data_flow = n6237_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:377:8  */
  assign wr_sram_data_flow = n6238_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:378:8  */
  assign wr_ddr_data_flow = n6239_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:379:8  */
  assign wr_stream = n6240_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:382:8  */
  assign wr_stream_id = n6243_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:386:8  */
  assign log1 = dp_gen_core_i_n5207; // (signal)
  /* ../../HW/src/dp/dp.vhd:387:8  */
  assign log1_valid = dp_gen_core_i_n5208; // (signal)
  /* ../../HW/src/dp/dp.vhd:388:8  */
  assign log2 = dp_gen_core_i_n5209; // (signal)
  /* ../../HW/src/dp/dp.vhd:389:8  */
  assign log2_valid = dp_gen_core_i_n5210; // (signal)
  /* ../../HW/src/dp/dp.vhd:391:8  */
  assign readmaster1_addr = dp_source1_i_n5534; // (signal)
  /* ../../HW/src/dp/dp.vhd:392:8  */
  assign readmaster2_addr = dp_source2_i_n5686; // (signal)
  /* ../../HW/src/dp/dp.vhd:393:8  */
  assign readmaster3_addr = dp_source3_i0_n5832; // (signal)
  /* ../../HW/src/dp/dp.vhd:394:8  */
  assign writemaster1_addr = dp_sink1_i_n5979; // (signal)
  /* ../../HW/src/dp/dp.vhd:395:8  */
  assign writemaster2_addr = dp_sink2_i_n6051; // (signal)
  /* ../../HW/src/dp/dp.vhd:396:8  */
  assign writemaster3_addr = dp_sink3_i_n6118; // (signal)
  /* ../../HW/src/dp/dp.vhd:400:61  */
  assign n5147_o = readmaster1_addr[21:0];
  /* ../../HW/src/dp/dp.vhd:401:61  */
  assign n5148_o = readmaster2_addr[17:0];
  /* ../../HW/src/dp/dp.vhd:403:56  */
  assign n5149_o = wr_data[143:128];
  /* ../../HW/src/dp/dp.vhd:404:63  */
  assign n5150_o = writemaster1_addr[21:0];
  /* ../../HW/src/dp/dp.vhd:405:63  */
  assign n5151_o = writemaster2_addr[17:0];
  /* ../../HW/src/dp/dp.vhd:439:47  */
  assign dp_fetch_1_i_n5153 = dp_fetch_1_i_bus_readdata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:440:52  */
  assign dp_fetch_1_i_n5154 = dp_fetch_1_i_bus_readdatavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:441:48  */
  assign dp_fetch_1_i_n5155 = dp_fetch_1_i_bus_writewait_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:442:47  */
  assign dp_fetch_1_i_n5156 = dp_fetch_1_i_bus_readwait_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:444:52  */
  assign dp_fetch_1_i_n5157 = dp_fetch_1_i_instruction_valid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:445:46  */
  assign dp_fetch_1_i_n5158 = n5175_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:446:50  */
  assign dp_fetch_1_i_n5159 = n5177_o; // (signal)
  /* ../../HW/src/dp/dp.vhd:452:52  */
  assign dp_fetch_1_i_n5160 = dp_fetch_1_i_task_start_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:454:49  */
  assign dp_fetch_1_i_n5161 = dp_fetch_1_i_task_pending_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:453:41  */
  assign dp_fetch_1_i_n5162 = dp_fetch_1_i_task_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:455:44  */
  assign dp_fetch_1_i_n5163 = dp_fetch_1_i_task_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:456:46  */
  assign dp_fetch_1_i_n5164 = dp_fetch_1_i_task_pcore_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:457:50  */
  assign dp_fetch_1_i_n5165 = dp_fetch_1_i_task_lockstep_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:458:50  */
  assign dp_fetch_1_i_n5166 = dp_fetch_1_i_task_tid_mask_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:459:56  */
  assign dp_fetch_1_i_n5167 = dp_fetch_1_i_task_iregister_auto_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:460:52  */
  assign dp_fetch_1_i_n5168 = dp_fetch_1_i_task_data_model_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:464:53  */
  assign dp_fetch_1_i_n5169 = dp_fetch_1_i_indication_avail_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:425:1  */
  dp_fetch_0_3_3 dp_fetch_1_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .bus_waddr_in(bus_waddr_in),
    .bus_raddr_in(bus_raddr_in),
    .bus_write_in(bus_write_in),
    .bus_read_in(bus_read_in),
    .bus_writedata_in(bus_writedata_in),
    .ready_in(ready),
    .pcore_sink_counter_in(writemaster1_counter_in),
    .sram_sink_counter_in(writemaster2_counter_in),
    .ddr_sink_counter_in(writemaster3_counter_in),
    .task_busy_in(task_busy_in),
    .task_ready_in(task_ready_in),
    .log1_in(log1),
    .log1_valid_in(log1_valid),
    .log2_in(log2),
    .log2_valid_in(log2_valid),
    .pcore_read_pending_p0_in(pcore_read_pending_p0),
    .sram_read_pending_p0_in(sram_read_pending_p0),
    .ddr_read_pending_p0_in(ddr_read_pending_p0),
    .pcore_read_pending_p1_in(pcore_read_pending_p1),
    .sram_read_pending_p1_in(sram_read_pending_p1),
    .ddr_read_pending_p1_in(ddr_read_pending_p1),
    .ddr_tx_busy_in(ddr_tx_busy_in),
    .bus_readdata_out(dp_fetch_1_i_bus_readdata_out),
    .bus_readdatavalid_out(dp_fetch_1_i_bus_readdatavalid_out),
    .bus_writewait_out(dp_fetch_1_i_bus_writewait_out),
    .bus_readwait_out(dp_fetch_1_i_bus_readwait_out),
    .instruction_valid_out(dp_fetch_1_i_instruction_valid_out),
    .instruction_out_opcode(dp_fetch_1_i_instruction_out_opcode),
    .instruction_out_condition(dp_fetch_1_i_instruction_out_condition),
    .instruction_out_vm(dp_fetch_1_i_instruction_out_vm),
    .instruction_out_source(dp_fetch_1_i_instruction_out_source),
    .instruction_out_source_bus_id(dp_fetch_1_i_instruction_out_source_bus_id),
    .instruction_out_source_data_type(dp_fetch_1_i_instruction_out_source_data_type),
    .instruction_out_dest(dp_fetch_1_i_instruction_out_dest),
    .instruction_out_dest_bus_id(dp_fetch_1_i_instruction_out_dest_bus_id),
    .instruction_out_dest_data_type(dp_fetch_1_i_instruction_out_dest_data_type),
    .instruction_out_mcast(dp_fetch_1_i_instruction_out_mcast),
    .instruction_out_count(dp_fetch_1_i_instruction_out_count),
    .instruction_out_data(dp_fetch_1_i_instruction_out_data),
    .instruction_out_repeat(dp_fetch_1_i_instruction_out_repeat),
    .instruction_out_source_addr_mode(dp_fetch_1_i_instruction_out_source_addr_mode),
    .instruction_out_dest_addr_mode(dp_fetch_1_i_instruction_out_dest_addr_mode),
    .instruction_out_stream_process(dp_fetch_1_i_instruction_out_stream_process),
    .instruction_out_stream_process_id(dp_fetch_1_i_instruction_out_stream_process_id),
    .pre_instruction_out_opcode(dp_fetch_1_i_pre_instruction_out_opcode),
    .pre_instruction_out_condition(dp_fetch_1_i_pre_instruction_out_condition),
    .pre_instruction_out_vm(dp_fetch_1_i_pre_instruction_out_vm),
    .pre_instruction_out_source(dp_fetch_1_i_pre_instruction_out_source),
    .pre_instruction_out_source_bus_id(dp_fetch_1_i_pre_instruction_out_source_bus_id),
    .pre_instruction_out_source_data_type(dp_fetch_1_i_pre_instruction_out_source_data_type),
    .pre_instruction_out_dest(dp_fetch_1_i_pre_instruction_out_dest),
    .pre_instruction_out_dest_bus_id(dp_fetch_1_i_pre_instruction_out_dest_bus_id),
    .pre_instruction_out_dest_data_type(dp_fetch_1_i_pre_instruction_out_dest_data_type),
    .pre_instruction_out_mcast(dp_fetch_1_i_pre_instruction_out_mcast),
    .pre_instruction_out_count(dp_fetch_1_i_pre_instruction_out_count),
    .pre_instruction_out_data(dp_fetch_1_i_pre_instruction_out_data),
    .pre_instruction_out_repeat(dp_fetch_1_i_pre_instruction_out_repeat),
    .pre_instruction_out_source_addr_mode(dp_fetch_1_i_pre_instruction_out_source_addr_mode),
    .pre_instruction_out_dest_addr_mode(dp_fetch_1_i_pre_instruction_out_dest_addr_mode),
    .pre_instruction_out_stream_process(dp_fetch_1_i_pre_instruction_out_stream_process),
    .pre_instruction_out_stream_process_id(dp_fetch_1_i_pre_instruction_out_stream_process_id),
    .task_start_addr_out(dp_fetch_1_i_task_start_addr_out),
    .task_pending_out(dp_fetch_1_i_task_pending_out),
    .task_out(dp_fetch_1_i_task_out),
    .task_vm_out(dp_fetch_1_i_task_vm_out),
    .task_pcore_out(dp_fetch_1_i_task_pcore_out),
    .task_lockstep_out(dp_fetch_1_i_task_lockstep_out),
    .task_tid_mask_out(dp_fetch_1_i_task_tid_mask_out),
    .task_iregister_auto_out(dp_fetch_1_i_task_iregister_auto_out),
    .task_data_model_out(dp_fetch_1_i_task_data_model_out),
    .indication_avail_out(dp_fetch_1_i_indication_avail_out));
  assign n5175_o = {dp_fetch_1_i_instruction_out_stream_process_id, dp_fetch_1_i_instruction_out_stream_process, dp_fetch_1_i_instruction_out_dest_addr_mode, dp_fetch_1_i_instruction_out_source_addr_mode, dp_fetch_1_i_instruction_out_repeat, dp_fetch_1_i_instruction_out_data, dp_fetch_1_i_instruction_out_count, dp_fetch_1_i_instruction_out_mcast, dp_fetch_1_i_instruction_out_dest_data_type, dp_fetch_1_i_instruction_out_dest_bus_id, dp_fetch_1_i_instruction_out_dest, dp_fetch_1_i_instruction_out_source_data_type, dp_fetch_1_i_instruction_out_source_bus_id, dp_fetch_1_i_instruction_out_source, dp_fetch_1_i_instruction_out_vm, dp_fetch_1_i_instruction_out_condition, dp_fetch_1_i_instruction_out_opcode};
  assign n5177_o = {dp_fetch_1_i_pre_instruction_out_stream_process_id, dp_fetch_1_i_pre_instruction_out_stream_process, dp_fetch_1_i_pre_instruction_out_dest_addr_mode, dp_fetch_1_i_pre_instruction_out_source_addr_mode, dp_fetch_1_i_pre_instruction_out_repeat, dp_fetch_1_i_pre_instruction_out_data, dp_fetch_1_i_pre_instruction_out_count, dp_fetch_1_i_pre_instruction_out_mcast, dp_fetch_1_i_pre_instruction_out_dest_data_type, dp_fetch_1_i_pre_instruction_out_dest_bus_id, dp_fetch_1_i_pre_instruction_out_dest, dp_fetch_1_i_pre_instruction_out_source_data_type, dp_fetch_1_i_pre_instruction_out_source_bus_id, dp_fetch_1_i_pre_instruction_out_source, dp_fetch_1_i_pre_instruction_out_vm, dp_fetch_1_i_pre_instruction_out_condition, dp_fetch_1_i_pre_instruction_out_opcode};
  /* ../../HW/src/dp/dp.vhd:490:19  */
  assign dp_gen_core_i_n5206 = dp_gen_core_i_ready_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:499:18  */
  assign dp_gen_core_i_n5207 = dp_gen_core_i_log1_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:500:24  */
  assign dp_gen_core_i_n5208 = dp_gen_core_i_log1_valid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:502:18  */
  assign dp_gen_core_i_n5209 = dp_gen_core_i_log2_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:503:24  */
  assign dp_gen_core_i_n5210 = dp_gen_core_i_log2_valid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:507:34  */
  assign dp_gen_core_i_n5211 = dp_gen_core_i_gen_pcore_src_valid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:508:28  */
  assign dp_gen_core_i_n5212 = dp_gen_core_i_gen_pcore_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:509:29  */
  assign dp_gen_core_i_n5213 = dp_gen_core_i_gen_pcore_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:510:34  */
  assign dp_gen_core_i_n5214 = dp_gen_core_i_gen_pcore_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:511:35  */
  assign dp_gen_core_i_n5215 = dp_gen_core_i_gen_pcore_src_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:512:36  */
  assign dp_gen_core_i_n5216 = dp_gen_core_i_gen_pcore_dest_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:513:34  */
  assign dp_gen_core_i_n5217 = dp_gen_core_i_gen_pcore_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:514:35  */
  assign dp_gen_core_i_n5218 = dp_gen_core_i_gen_pcore_src_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:515:35  */
  assign dp_gen_core_i_n5219 = dp_gen_core_i_gen_pcore_dst_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:516:36  */
  assign dp_gen_core_i_n5220 = dp_gen_core_i_gen_pcore_src_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:517:36  */
  assign dp_gen_core_i_n5221 = dp_gen_core_i_gen_pcore_dst_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:518:34  */
  assign dp_gen_core_i_n5222 = dp_gen_core_i_gen_pcore_src_start_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:519:32  */
  assign dp_gen_core_i_n5223 = dp_gen_core_i_gen_pcore_src_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:520:32  */
  assign dp_gen_core_i_n5224 = dp_gen_core_i_gen_pcore_dst_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:521:33  */
  assign dp_gen_core_i_n5225 = dp_gen_core_i_gen_pcore_src_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:522:38  */
  assign dp_gen_core_i_n5226 = dp_gen_core_i_gen_pcore_src_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:523:33  */
  assign dp_gen_core_i_n5227 = dp_gen_core_i_gen_pcore_dst_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:524:38  */
  assign dp_gen_core_i_n5228 = dp_gen_core_i_gen_pcore_dst_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:525:32  */
  assign dp_gen_core_i_n5229 = dp_gen_core_i_gen_pcore_src_eof_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:526:38  */
  assign dp_gen_core_i_n5230 = dp_gen_core_i_gen_pcore_bus_id_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:527:41  */
  assign dp_gen_core_i_n5231 = dp_gen_core_i_gen_pcore_data_type_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:528:42  */
  assign dp_gen_core_i_n5232 = dp_gen_core_i_gen_pcore_data_model_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:529:36  */
  assign dp_gen_core_i_n5233 = dp_gen_core_i_gen_pcore_bus_id_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:530:34  */
  assign dp_gen_core_i_n5234 = dp_gen_core_i_gen_pcore_busy_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:531:39  */
  assign dp_gen_core_i_n5235 = dp_gen_core_i_gen_pcore_data_type_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:532:40  */
  assign dp_gen_core_i_n5236 = dp_gen_core_i_gen_pcore_data_model_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:533:37  */
  assign dp_gen_core_i_n5237 = dp_gen_core_i_gen_pcore_src_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:534:37  */
  assign dp_gen_core_i_n5238 = dp_gen_core_i_gen_pcore_dst_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:535:31  */
  assign dp_gen_core_i_n5239 = dp_gen_core_i_gen_pcore_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:536:30  */
  assign dp_gen_core_i_n5240 = dp_gen_core_i_gen_pcore_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:537:29  */
  assign dp_gen_core_i_n5241 = dp_gen_core_i_gen_pcore_data_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:541:33  */
  assign dp_gen_core_i_n5242 = dp_gen_core_i_gen_sram_src_valid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:542:27  */
  assign dp_gen_core_i_n5243 = dp_gen_core_i_gen_sram_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:543:28  */
  assign dp_gen_core_i_n5244 = dp_gen_core_i_gen_sram_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:544:33  */
  assign dp_gen_core_i_n5245 = dp_gen_core_i_gen_sram_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:545:34  */
  assign dp_gen_core_i_n5246 = dp_gen_core_i_gen_sram_src_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:546:35  */
  assign dp_gen_core_i_n5247 = dp_gen_core_i_gen_sram_dest_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:547:33  */
  assign dp_gen_core_i_n5248 = dp_gen_core_i_gen_sram_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:548:34  */
  assign dp_gen_core_i_n5249 = dp_gen_core_i_gen_sram_src_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:549:34  */
  assign dp_gen_core_i_n5250 = dp_gen_core_i_gen_sram_dst_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:550:35  */
  assign dp_gen_core_i_n5251 = dp_gen_core_i_gen_sram_src_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:551:35  */
  assign dp_gen_core_i_n5252 = dp_gen_core_i_gen_sram_dst_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:552:33  */
  assign dp_gen_core_i_n5253 = dp_gen_core_i_gen_sram_src_start_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:553:31  */
  assign dp_gen_core_i_n5254 = dp_gen_core_i_gen_sram_src_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:554:31  */
  assign dp_gen_core_i_n5255 = dp_gen_core_i_gen_sram_dst_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:555:32  */
  assign dp_gen_core_i_n5256 = dp_gen_core_i_gen_sram_src_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:556:37  */
  assign dp_gen_core_i_n5257 = dp_gen_core_i_gen_sram_src_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:557:32  */
  assign dp_gen_core_i_n5258 = dp_gen_core_i_gen_sram_dst_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:558:37  */
  assign dp_gen_core_i_n5259 = dp_gen_core_i_gen_sram_dst_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:559:31  */
  assign dp_gen_core_i_n5260 = dp_gen_core_i_gen_sram_src_eof_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:560:37  */
  assign dp_gen_core_i_n5261 = dp_gen_core_i_gen_sram_bus_id_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:561:40  */
  assign dp_gen_core_i_n5262 = dp_gen_core_i_gen_sram_data_type_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:562:41  */
  assign dp_gen_core_i_n5263 = dp_gen_core_i_gen_sram_data_model_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:563:35  */
  assign dp_gen_core_i_n5264 = dp_gen_core_i_gen_sram_bus_id_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:564:33  */
  assign dp_gen_core_i_n5265 = dp_gen_core_i_gen_sram_busy_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:565:38  */
  assign dp_gen_core_i_n5266 = dp_gen_core_i_gen_sram_data_type_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:566:39  */
  assign dp_gen_core_i_n5267 = dp_gen_core_i_gen_sram_data_model_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:567:36  */
  assign dp_gen_core_i_n5268 = dp_gen_core_i_gen_sram_src_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:568:36  */
  assign dp_gen_core_i_n5269 = dp_gen_core_i_gen_sram_dst_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:569:30  */
  assign dp_gen_core_i_n5270 = dp_gen_core_i_gen_sram_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:570:29  */
  assign dp_gen_core_i_n5271 = dp_gen_core_i_gen_sram_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:571:28  */
  assign dp_gen_core_i_n5272 = dp_gen_core_i_gen_sram_data_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:575:32  */
  assign dp_gen_core_i_n5273 = dp_gen_core_i_gen_ddr_src_valid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:576:26  */
  assign dp_gen_core_i_n5274 = dp_gen_core_i_gen_ddr_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:577:27  */
  assign dp_gen_core_i_n5275 = dp_gen_core_i_gen_ddr_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:578:32  */
  assign dp_gen_core_i_n5276 = dp_gen_core_i_gen_ddr_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:579:33  */
  assign dp_gen_core_i_n5277 = dp_gen_core_i_gen_ddr_src_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:580:34  */
  assign dp_gen_core_i_n5278 = dp_gen_core_i_gen_ddr_dest_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:581:32  */
  assign dp_gen_core_i_n5279 = dp_gen_core_i_gen_ddr_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:582:33  */
  assign dp_gen_core_i_n5280 = dp_gen_core_i_gen_ddr_src_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:583:33  */
  assign dp_gen_core_i_n5281 = dp_gen_core_i_gen_ddr_dst_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:584:34  */
  assign dp_gen_core_i_n5282 = dp_gen_core_i_gen_ddr_src_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:585:34  */
  assign dp_gen_core_i_n5283 = dp_gen_core_i_gen_ddr_dst_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:586:32  */
  assign dp_gen_core_i_n5284 = dp_gen_core_i_gen_ddr_src_start_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:587:30  */
  assign dp_gen_core_i_n5285 = dp_gen_core_i_gen_ddr_src_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:588:30  */
  assign dp_gen_core_i_n5286 = dp_gen_core_i_gen_ddr_dst_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:589:31  */
  assign dp_gen_core_i_n5287 = dp_gen_core_i_gen_ddr_src_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:590:36  */
  assign dp_gen_core_i_n5288 = dp_gen_core_i_gen_ddr_src_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:591:31  */
  assign dp_gen_core_i_n5289 = dp_gen_core_i_gen_ddr_dst_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:592:36  */
  assign dp_gen_core_i_n5290 = dp_gen_core_i_gen_ddr_dst_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:593:30  */
  assign dp_gen_core_i_n5291 = dp_gen_core_i_gen_ddr_src_eof_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:594:36  */
  assign dp_gen_core_i_n5292 = dp_gen_core_i_gen_ddr_bus_id_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:595:39  */
  assign dp_gen_core_i_n5293 = dp_gen_core_i_gen_ddr_data_type_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:596:40  */
  assign dp_gen_core_i_n5294 = dp_gen_core_i_gen_ddr_data_model_source_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:597:34  */
  assign dp_gen_core_i_n5295 = dp_gen_core_i_gen_ddr_bus_id_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:598:32  */
  assign dp_gen_core_i_n5296 = dp_gen_core_i_gen_ddr_busy_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:599:37  */
  assign dp_gen_core_i_n5297 = dp_gen_core_i_gen_ddr_data_type_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:600:38  */
  assign dp_gen_core_i_n5298 = dp_gen_core_i_gen_ddr_data_model_dest_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:601:35  */
  assign dp_gen_core_i_n5299 = dp_gen_core_i_gen_ddr_src_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:602:35  */
  assign dp_gen_core_i_n5300 = dp_gen_core_i_gen_ddr_dst_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:603:29  */
  assign dp_gen_core_i_n5301 = dp_gen_core_i_gen_ddr_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:604:28  */
  assign dp_gen_core_i_n5302 = dp_gen_core_i_gen_ddr_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:605:27  */
  assign dp_gen_core_i_n5303 = dp_gen_core_i_gen_ddr_data_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:483:1  */
  dp_gen_core dp_gen_core_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .instruction_valid_in(valid),
    .instruction_in_opcode(n5305_o),
    .instruction_in_condition(n5306_o),
    .instruction_in_vm(n5307_o),
    .instruction_in_source(n5308_o),
    .instruction_in_source_bus_id(n5309_o),
    .instruction_in_source_data_type(n5310_o),
    .instruction_in_dest(n5311_o),
    .instruction_in_dest_bus_id(n5312_o),
    .instruction_in_dest_data_type(n5313_o),
    .instruction_in_mcast(n5314_o),
    .instruction_in_count(n5315_o),
    .instruction_in_data(n5316_o),
    .instruction_in_repeat(n5317_o),
    .instruction_in_source_addr_mode(n5318_o),
    .instruction_in_dest_addr_mode(n5319_o),
    .instruction_in_stream_process(n5320_o),
    .instruction_in_stream_process_id(n5321_o),
    .pre_instruction_in_opcode(n5322_o),
    .pre_instruction_in_condition(n5323_o),
    .pre_instruction_in_vm(n5324_o),
    .pre_instruction_in_source(n5325_o),
    .pre_instruction_in_source_bus_id(n5326_o),
    .pre_instruction_in_source_data_type(n5327_o),
    .pre_instruction_in_dest(n5328_o),
    .pre_instruction_in_dest_bus_id(n5329_o),
    .pre_instruction_in_dest_data_type(n5330_o),
    .pre_instruction_in_mcast(n5331_o),
    .pre_instruction_in_count(n5332_o),
    .pre_instruction_in_data(n5333_o),
    .pre_instruction_in_repeat(n5334_o),
    .pre_instruction_in_source_addr_mode(n5335_o),
    .pre_instruction_in_dest_addr_mode(n5336_o),
    .pre_instruction_in_stream_process(n5337_o),
    .pre_instruction_in_stream_process_id(n5338_o),
    .wr_maxburstlen_in(wr_maxburstlen),
    .full_in(full),
    .waitreq_in(waitreq),
    .bar_in(bar_in),
    .ready_out(dp_gen_core_i_ready_out),
    .log1_out(dp_gen_core_i_log1_out),
    .log1_valid_out(dp_gen_core_i_log1_valid_out),
    .log2_out(dp_gen_core_i_log2_out),
    .log2_valid_out(dp_gen_core_i_log2_valid_out),
    .gen_pcore_src_valid_out(dp_gen_core_i_gen_pcore_src_valid_out),
    .gen_pcore_vm_out(dp_gen_core_i_gen_pcore_vm_out),
    .gen_pcore_fork_out(dp_gen_core_i_gen_pcore_fork_out),
    .gen_pcore_data_flow_out(dp_gen_core_i_gen_pcore_data_flow_out),
    .gen_pcore_src_stream_out(dp_gen_core_i_gen_pcore_src_stream_out),
    .gen_pcore_dest_stream_out(dp_gen_core_i_gen_pcore_dest_stream_out),
    .gen_pcore_stream_id_out(dp_gen_core_i_gen_pcore_stream_id_out),
    .gen_pcore_src_vector_out(dp_gen_core_i_gen_pcore_src_vector_out),
    .gen_pcore_dst_vector_out(dp_gen_core_i_gen_pcore_dst_vector_out),
    .gen_pcore_src_scatter_out(dp_gen_core_i_gen_pcore_src_scatter_out),
    .gen_pcore_dst_scatter_out(dp_gen_core_i_gen_pcore_dst_scatter_out),
    .gen_pcore_src_start_out(dp_gen_core_i_gen_pcore_src_start_out),
    .gen_pcore_src_end_out(dp_gen_core_i_gen_pcore_src_end_out),
    .gen_pcore_dst_end_out(dp_gen_core_i_gen_pcore_dst_end_out),
    .gen_pcore_src_addr_out(dp_gen_core_i_gen_pcore_src_addr_out),
    .gen_pcore_src_addr_mode_out(dp_gen_core_i_gen_pcore_src_addr_mode_out),
    .gen_pcore_dst_addr_out(dp_gen_core_i_gen_pcore_dst_addr_out),
    .gen_pcore_dst_addr_mode_out(dp_gen_core_i_gen_pcore_dst_addr_mode_out),
    .gen_pcore_src_eof_out(dp_gen_core_i_gen_pcore_src_eof_out),
    .gen_pcore_bus_id_source_out(dp_gen_core_i_gen_pcore_bus_id_source_out),
    .gen_pcore_data_type_source_out(dp_gen_core_i_gen_pcore_data_type_source_out),
    .gen_pcore_data_model_source_out(dp_gen_core_i_gen_pcore_data_model_source_out),
    .gen_pcore_bus_id_dest_out(dp_gen_core_i_gen_pcore_bus_id_dest_out),
    .gen_pcore_busy_dest_out(dp_gen_core_i_gen_pcore_busy_dest_out),
    .gen_pcore_data_type_dest_out(dp_gen_core_i_gen_pcore_data_type_dest_out),
    .gen_pcore_data_model_dest_out(dp_gen_core_i_gen_pcore_data_model_dest_out),
    .gen_pcore_src_burstlen_out(dp_gen_core_i_gen_pcore_src_burstlen_out),
    .gen_pcore_dst_burstlen_out(dp_gen_core_i_gen_pcore_dst_burstlen_out),
    .gen_pcore_thread_out(dp_gen_core_i_gen_pcore_thread_out),
    .gen_pcore_mcast_out(dp_gen_core_i_gen_pcore_mcast_out),
    .gen_pcore_data_out(dp_gen_core_i_gen_pcore_data_out),
    .gen_sram_src_valid_out(dp_gen_core_i_gen_sram_src_valid_out),
    .gen_sram_vm_out(dp_gen_core_i_gen_sram_vm_out),
    .gen_sram_fork_out(dp_gen_core_i_gen_sram_fork_out),
    .gen_sram_data_flow_out(dp_gen_core_i_gen_sram_data_flow_out),
    .gen_sram_src_stream_out(dp_gen_core_i_gen_sram_src_stream_out),
    .gen_sram_dest_stream_out(dp_gen_core_i_gen_sram_dest_stream_out),
    .gen_sram_stream_id_out(dp_gen_core_i_gen_sram_stream_id_out),
    .gen_sram_src_vector_out(dp_gen_core_i_gen_sram_src_vector_out),
    .gen_sram_dst_vector_out(dp_gen_core_i_gen_sram_dst_vector_out),
    .gen_sram_src_scatter_out(dp_gen_core_i_gen_sram_src_scatter_out),
    .gen_sram_dst_scatter_out(dp_gen_core_i_gen_sram_dst_scatter_out),
    .gen_sram_src_start_out(dp_gen_core_i_gen_sram_src_start_out),
    .gen_sram_src_end_out(dp_gen_core_i_gen_sram_src_end_out),
    .gen_sram_dst_end_out(dp_gen_core_i_gen_sram_dst_end_out),
    .gen_sram_src_addr_out(dp_gen_core_i_gen_sram_src_addr_out),
    .gen_sram_src_addr_mode_out(dp_gen_core_i_gen_sram_src_addr_mode_out),
    .gen_sram_dst_addr_out(dp_gen_core_i_gen_sram_dst_addr_out),
    .gen_sram_dst_addr_mode_out(dp_gen_core_i_gen_sram_dst_addr_mode_out),
    .gen_sram_src_eof_out(dp_gen_core_i_gen_sram_src_eof_out),
    .gen_sram_bus_id_source_out(dp_gen_core_i_gen_sram_bus_id_source_out),
    .gen_sram_data_type_source_out(dp_gen_core_i_gen_sram_data_type_source_out),
    .gen_sram_data_model_source_out(dp_gen_core_i_gen_sram_data_model_source_out),
    .gen_sram_bus_id_dest_out(dp_gen_core_i_gen_sram_bus_id_dest_out),
    .gen_sram_busy_dest_out(dp_gen_core_i_gen_sram_busy_dest_out),
    .gen_sram_data_type_dest_out(dp_gen_core_i_gen_sram_data_type_dest_out),
    .gen_sram_data_model_dest_out(dp_gen_core_i_gen_sram_data_model_dest_out),
    .gen_sram_src_burstlen_out(dp_gen_core_i_gen_sram_src_burstlen_out),
    .gen_sram_dst_burstlen_out(dp_gen_core_i_gen_sram_dst_burstlen_out),
    .gen_sram_thread_out(dp_gen_core_i_gen_sram_thread_out),
    .gen_sram_mcast_out(dp_gen_core_i_gen_sram_mcast_out),
    .gen_sram_data_out(dp_gen_core_i_gen_sram_data_out),
    .gen_ddr_src_valid_out(dp_gen_core_i_gen_ddr_src_valid_out),
    .gen_ddr_vm_out(dp_gen_core_i_gen_ddr_vm_out),
    .gen_ddr_fork_out(dp_gen_core_i_gen_ddr_fork_out),
    .gen_ddr_data_flow_out(dp_gen_core_i_gen_ddr_data_flow_out),
    .gen_ddr_src_stream_out(dp_gen_core_i_gen_ddr_src_stream_out),
    .gen_ddr_dest_stream_out(dp_gen_core_i_gen_ddr_dest_stream_out),
    .gen_ddr_stream_id_out(dp_gen_core_i_gen_ddr_stream_id_out),
    .gen_ddr_src_vector_out(dp_gen_core_i_gen_ddr_src_vector_out),
    .gen_ddr_dst_vector_out(dp_gen_core_i_gen_ddr_dst_vector_out),
    .gen_ddr_src_scatter_out(dp_gen_core_i_gen_ddr_src_scatter_out),
    .gen_ddr_dst_scatter_out(dp_gen_core_i_gen_ddr_dst_scatter_out),
    .gen_ddr_src_start_out(dp_gen_core_i_gen_ddr_src_start_out),
    .gen_ddr_src_end_out(dp_gen_core_i_gen_ddr_src_end_out),
    .gen_ddr_dst_end_out(dp_gen_core_i_gen_ddr_dst_end_out),
    .gen_ddr_src_addr_out(dp_gen_core_i_gen_ddr_src_addr_out),
    .gen_ddr_src_addr_mode_out(dp_gen_core_i_gen_ddr_src_addr_mode_out),
    .gen_ddr_dst_addr_out(dp_gen_core_i_gen_ddr_dst_addr_out),
    .gen_ddr_dst_addr_mode_out(dp_gen_core_i_gen_ddr_dst_addr_mode_out),
    .gen_ddr_src_eof_out(dp_gen_core_i_gen_ddr_src_eof_out),
    .gen_ddr_bus_id_source_out(dp_gen_core_i_gen_ddr_bus_id_source_out),
    .gen_ddr_data_type_source_out(dp_gen_core_i_gen_ddr_data_type_source_out),
    .gen_ddr_data_model_source_out(dp_gen_core_i_gen_ddr_data_model_source_out),
    .gen_ddr_bus_id_dest_out(dp_gen_core_i_gen_ddr_bus_id_dest_out),
    .gen_ddr_busy_dest_out(dp_gen_core_i_gen_ddr_busy_dest_out),
    .gen_ddr_data_type_dest_out(dp_gen_core_i_gen_ddr_data_type_dest_out),
    .gen_ddr_data_model_dest_out(dp_gen_core_i_gen_ddr_data_model_dest_out),
    .gen_ddr_src_burstlen_out(dp_gen_core_i_gen_ddr_src_burstlen_out),
    .gen_ddr_dst_burstlen_out(dp_gen_core_i_gen_ddr_dst_burstlen_out),
    .gen_ddr_thread_out(dp_gen_core_i_gen_ddr_thread_out),
    .gen_ddr_mcast_out(dp_gen_core_i_gen_ddr_mcast_out),
    .gen_ddr_data_out(dp_gen_core_i_gen_ddr_data_out));
  assign n5305_o = instruction[2:0];
  assign n5306_o = instruction[6:3];
  assign n5307_o = instruction[7];
  assign n5308_o = instruction[783:8];
  assign n5309_o = instruction[785:784];
  assign n5310_o = instruction[787:786];
  assign n5311_o = instruction[1563:788];
  assign n5312_o = instruction[1565:1564];
  assign n5313_o = instruction[1567:1566];
  assign n5314_o = instruction[1573:1568];
  assign n5315_o = instruction[1597:1574];
  assign n5316_o = instruction[1613:1598];
  assign n5317_o = instruction[1614];
  assign n5318_o = instruction[1615];
  assign n5319_o = instruction[1616];
  assign n5320_o = instruction[1617];
  assign n5321_o = instruction[1619:1618];
  assign n5322_o = pre_instruction[2:0];
  assign n5323_o = pre_instruction[6:3];
  assign n5324_o = pre_instruction[7];
  assign n5325_o = pre_instruction[783:8];
  assign n5326_o = pre_instruction[785:784];
  assign n5327_o = pre_instruction[787:786];
  assign n5328_o = pre_instruction[1563:788];
  assign n5329_o = pre_instruction[1565:1564];
  assign n5330_o = pre_instruction[1567:1566];
  assign n5331_o = pre_instruction[1573:1568];
  assign n5332_o = pre_instruction[1597:1574];
  assign n5333_o = pre_instruction[1613:1598];
  assign n5334_o = pre_instruction[1614];
  assign n5335_o = pre_instruction[1615];
  assign n5336_o = pre_instruction[1616];
  assign n5337_o = pre_instruction[1617];
  assign n5338_o = pre_instruction[1619:1618];
  /* ../../HW/src/dp/dp.vhd:625:27  */
  assign dp_source1_i_n5534 = dp_source1_i_bus_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:626:32  */
  assign dp_source1_i_n5535 = dp_source1_i_bus_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:627:25  */
  assign dp_source1_i_n5536 = dp_source1_i_bus_cs_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:628:27  */
  assign dp_source1_i_n5537 = dp_source1_i_bus_read_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:629:30  */
  assign dp_source1_i_n5538 = dp_source1_i_bus_read_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:630:32  */
  assign dp_source1_i_n5539 = dp_source1_i_bus_read_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:631:37  */
  assign dp_source1_i_n5540 = dp_source1_i_bus_read_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:632:34  */
  assign dp_source1_i_n5541 = dp_source1_i_bus_read_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:633:37  */
  assign dp_source1_i_n5542 = dp_source1_i_bus_read_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:634:34  */
  assign dp_source1_i_n5543 = dp_source1_i_bus_read_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:635:35  */
  assign dp_source1_i_n5544 = dp_source1_i_bus_read_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:642:31  */
  assign dp_source1_i_n5547 = dp_source1_i_bus_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:643:25  */
  assign dp_source1_i_n5548 = dp_source1_i_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:644:32  */
  assign dp_source1_i_n5549 = dp_source1_i_bus_data_type_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:645:33  */
  assign dp_source1_i_n5550 = dp_source1_i_bus_data_model_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:647:30  */
  assign dp_source1_i_n5551 = dp_source1_i_gen_waitreq_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:680:29  */
  assign dp_source1_i_n5552 = dp_source1_i_wr_req_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:684:40  */
  assign dp_source1_i_n5553 = dp_source1_i_wr_req_pending_p0_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:688:40  */
  assign dp_source1_i_n5554 = dp_source1_i_wr_req_pending_p1_out; // (signal)
  assign n5555_o = {wr_ddr_full, wr_sram_full, wr_full};
  /* ../../HW/src/dp/dp.vhd:696:34  */
  assign dp_source1_i_n5556 = dp_source1_i_wr_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:700:31  */
  assign dp_source1_i_n5557 = dp_source1_i_wr_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:704:31  */
  assign dp_source1_i_n5558 = dp_source1_i_wr_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:708:34  */
  assign dp_source1_i_n5559 = dp_source1_i_wr_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:712:32  */
  assign dp_source1_i_n5560 = dp_source1_i_wr_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:716:28  */
  assign dp_source1_i_n5561 = dp_source1_i_wr_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:720:27  */
  assign dp_source1_i_n5562 = dp_source1_i_wr_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:722:27  */
  assign dp_source1_i_n5563 = dp_source1_i_wr_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:724:30  */
  assign dp_source1_i_n5564 = dp_source1_i_wr_src_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:726:31  */
  assign dp_source1_i_n5565 = dp_source1_i_wr_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:728:33  */
  assign dp_source1_i_n5566 = dp_source1_i_wr_datavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:730:27  */
  assign dp_source1_i_n5567 = dp_source1_i_wr_data_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:732:37  */
  assign dp_source1_i_n5568 = dp_source1_i_wr_readdatavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:734:40  */
  assign dp_source1_i_n5569 = dp_source1_i_wr_readdatavalid_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:736:32  */
  assign dp_source1_i_n5570 = dp_source1_i_wr_readdata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:738:31  */
  assign dp_source1_i_n5571 = dp_source1_i_wr_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:740:29  */
  assign dp_source1_i_n5572 = dp_source1_i_wr_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:742:28  */
  assign dp_source1_i_n5573 = dp_source1_i_wr_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:744:31  */
  assign dp_source1_i_n5574 = dp_source1_i_wr_data_type_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:746:32  */
  assign dp_source1_i_n5575 = dp_source1_i_wr_data_model_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:748:27  */
  assign dp_source1_i_n5576 = dp_source1_i_wr_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:612:1  */
  dp_source_0_3_8_32_1_0 dp_source1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .bus_readdatavalid_in(readmaster1_readdatavalid_in),
    .bus_readdatavalid_vm_in(readmaster1_readdatavalid_vm_in),
    .bus_readdata_in(readmaster1_readdata_in),
    .bus_wait_request_in(readmaster1_wait_request_in),
    .gen_valid_in(gen_pcore_src_valid),
    .gen_vm_in(gen_pcore_vm),
    .gen_fork_in(gen_pcore_fork),
    .gen_data_flow_in(gen_pcore_data_flow),
    .gen_src_stream_in(gen_pcore_src_stream),
    .gen_dest_stream_in(gen_pcore_dest_stream),
    .gen_stream_id_in(gen_pcore_stream_id),
    .gen_src_vector_in(gen_pcore_src_vector),
    .gen_dst_vector_in(gen_pcore_dst_vector),
    .gen_src_scatter_in(gen_pcore_src_scatter),
    .gen_dst_scatter_in(gen_pcore_dst_scatter),
    .gen_src_start_in(gen_pcore_src_start),
    .gen_src_end_in(gen_pcore_src_end),
    .gen_dst_end_in(gen_pcore_dst_end),
    .gen_src_eof_in(gen_pcore_src_eof),
    .gen_src_addr_in(gen_pcore_src_addr),
    .gen_src_addr_mode_in(gen_pcore_src_addr_mode),
    .gen_dst_addr_in(gen_pcore_dst_addr),
    .gen_dst_addr_mode_in(gen_pcore_dst_addr_mode),
    .gen_bus_id_source_in(gen_pcore_bus_id_source),
    .gen_data_type_source_in(gen_pcore_data_type_source),
    .gen_data_model_source_in(gen_pcore_data_model_source),
    .gen_bus_id_dest_in(gen_pcore_bus_id_dest),
    .gen_busy_dest_in(gen_pcore_busy_dest),
    .gen_data_type_dest_in(gen_pcore_data_type_dest),
    .gen_data_model_dest_in(gen_pcore_data_model_dest),
    .gen_src_burstlen_in(gen_pcore_src_burstlen),
    .gen_dst_burstlen_in(gen_pcore_dst_burstlen),
    .gen_thread_in(gen_pcore_thread),
    .gen_mcast_in(gen_pcore_mcast),
    .gen_src_data_in(gen_pcore_data),
    .wr_full_in(n5555_o),
    .bus_addr_out(dp_source1_i_bus_addr_out),
    .bus_addr_mode_out(dp_source1_i_bus_addr_mode_out),
    .bus_cs_out(dp_source1_i_bus_cs_out),
    .bus_read_out(dp_source1_i_bus_read_out),
    .bus_read_vm_out(dp_source1_i_bus_read_vm_out),
    .bus_read_fork_out(dp_source1_i_bus_read_fork_out),
    .bus_read_data_flow_out(dp_source1_i_bus_read_data_flow_out),
    .bus_read_stream_out(dp_source1_i_bus_read_stream_out),
    .bus_read_stream_id_out(dp_source1_i_bus_read_stream_id_out),
    .bus_read_vector_out(dp_source1_i_bus_read_vector_out),
    .bus_read_scatter_out(dp_source1_i_bus_read_scatter_out),
    .bus_read_start_out(),
    .bus_read_end_out(),
    .bus_burstlen_out(dp_source1_i_bus_burstlen_out),
    .bus_id_out(dp_source1_i_bus_id_out),
    .bus_data_type_out(dp_source1_i_bus_data_type_out),
    .bus_data_model_out(dp_source1_i_bus_data_model_out),
    .gen_waitreq_out(dp_source1_i_gen_waitreq_out),
    .wr_req_out(dp_source1_i_wr_req_out),
    .wr_req_pending_p0_out(dp_source1_i_wr_req_pending_p0_out),
    .wr_req_pending_p1_out(dp_source1_i_wr_req_pending_p1_out),
    .wr_data_flow_out(dp_source1_i_wr_data_flow_out),
    .wr_vector_out(dp_source1_i_wr_vector_out),
    .wr_stream_out(dp_source1_i_wr_stream_out),
    .wr_stream_id_out(dp_source1_i_wr_stream_id_out),
    .wr_scatter_out(dp_source1_i_wr_scatter_out),
    .wr_end_out(dp_source1_i_wr_end_out),
    .wr_addr_out(dp_source1_i_wr_addr_out),
    .wr_fork_out(dp_source1_i_wr_fork_out),
    .wr_addr_mode_out(dp_source1_i_wr_addr_mode_out),
    .wr_src_vm_out(dp_source1_i_wr_src_vm_out),
    .wr_datavalid_out(dp_source1_i_wr_datavalid_out),
    .wr_data_out(dp_source1_i_wr_data_out),
    .wr_readdatavalid_out(dp_source1_i_wr_readdatavalid_out),
    .wr_readdatavalid_vm_out(dp_source1_i_wr_readdatavalid_vm_out),
    .wr_readdata_out(dp_source1_i_wr_readdata_out),
    .wr_burstlen_out(dp_source1_i_wr_burstlen_out),
    .wr_bus_id_out(dp_source1_i_wr_bus_id_out),
    .wr_thread_out(dp_source1_i_wr_thread_out),
    .wr_data_type_out(dp_source1_i_wr_data_type_out),
    .wr_data_model_out(dp_source1_i_wr_data_model_out),
    .wr_mcast_out(dp_source1_i_wr_mcast_out));
  assign n5636_o = dp_source1_i_n5552[0];
  assign n5637_o = dp_source1_i_n5552[1];
  assign n5638_o = dp_source1_i_n5552[2];
  assign n5640_o = dp_source1_i_n5553[0];
  assign n5641_o = dp_source1_i_n5553[1];
  assign n5642_o = dp_source1_i_n5553[2];
  assign n5644_o = dp_source1_i_n5554[0];
  assign n5645_o = dp_source1_i_n5554[1];
  assign n5646_o = dp_source1_i_n5554[2];
  assign n5648_o = dp_source1_i_n5556[1:0];
  assign n5649_o = dp_source1_i_n5556[3:2];
  assign n5650_o = dp_source1_i_n5556[5:4];
  assign n5652_o = dp_source1_i_n5557[2:0];
  assign n5653_o = dp_source1_i_n5557[5:3];
  assign n5654_o = dp_source1_i_n5557[8:6];
  assign n5656_o = dp_source1_i_n5558[0];
  assign n5660_o = dp_source1_i_n5559[1:0];
  assign n5664_o = dp_source1_i_n5560[1:0];
  assign n5665_o = dp_source1_i_n5560[3:2];
  assign n5666_o = dp_source1_i_n5560[5:4];
  assign n5668_o = dp_source1_i_n5561[3:0];
  assign n5669_o = dp_source1_i_n5561[7:4];
  assign n5670_o = dp_source1_i_n5561[11:8];
  /* ../../HW/src/dp/dp.vhd:768:27  */
  assign dp_source2_i_n5686 = dp_source2_i_bus_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:769:25  */
  assign dp_source2_i_n5688 = dp_source2_i_bus_cs_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:770:27  */
  assign dp_source2_i_n5689 = dp_source2_i_bus_read_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:771:30  */
  assign dp_source2_i_n5690 = dp_source2_i_bus_read_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:772:32  */
  assign dp_source2_i_n5691 = dp_source2_i_bus_read_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:776:34  */
  assign dp_source2_i_n5695 = dp_source2_i_bus_read_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:777:35  */
  assign dp_source2_i_n5696 = dp_source2_i_bus_read_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:784:31  */
  assign dp_source2_i_n5699 = dp_source2_i_bus_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:785:25  */
  assign dp_source2_i_n5700 = dp_source2_i_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:789:30  */
  assign dp_source2_i_n5703 = dp_source2_i_gen_waitreq_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:822:29  */
  assign dp_source2_i_n5704 = dp_source2_i_wr_req_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:826:40  */
  assign dp_source2_i_n5705 = dp_source2_i_wr_req_pending_p0_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:830:40  */
  assign dp_source2_i_n5706 = dp_source2_i_wr_req_pending_p1_out; // (signal)
  assign n5707_o = {wr_ddr_full, wr_sram_full, wr_full};
  /* ../../HW/src/dp/dp.vhd:838:34  */
  assign dp_source2_i_n5708 = dp_source2_i_wr_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:842:31  */
  assign dp_source2_i_n5709 = dp_source2_i_wr_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:846:31  */
  assign dp_source2_i_n5710 = dp_source2_i_wr_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:850:34  */
  assign dp_source2_i_n5711 = dp_source2_i_wr_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:854:32  */
  assign dp_source2_i_n5712 = dp_source2_i_wr_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:858:28  */
  assign dp_source2_i_n5713 = dp_source2_i_wr_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:862:27  */
  assign dp_source2_i_n5714 = dp_source2_i_wr_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:864:27  */
  assign dp_source2_i_n5715 = dp_source2_i_wr_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:866:30  */
  assign dp_source2_i_n5716 = dp_source2_i_wr_src_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:868:31  */
  assign dp_source2_i_n5717 = dp_source2_i_wr_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:870:33  */
  assign dp_source2_i_n5718 = dp_source2_i_wr_datavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:872:27  */
  assign dp_source2_i_n5719 = dp_source2_i_wr_data_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:874:37  */
  assign dp_source2_i_n5720 = dp_source2_i_wr_readdatavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:876:40  */
  assign dp_source2_i_n5721 = dp_source2_i_wr_readdatavalid_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:878:32  */
  assign dp_source2_i_n5722 = dp_source2_i_wr_readdata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:880:31  */
  assign dp_source2_i_n5723 = dp_source2_i_wr_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:882:29  */
  assign dp_source2_i_n5724 = dp_source2_i_wr_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:884:28  */
  assign dp_source2_i_n5725 = dp_source2_i_wr_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:886:31  */
  assign dp_source2_i_n5726 = dp_source2_i_wr_data_type_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:888:32  */
  assign dp_source2_i_n5727 = dp_source2_i_wr_data_model_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:890:27  */
  assign dp_source2_i_n5728 = dp_source2_i_wr_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:755:1  */
  dp_source_1_3_4_32_1_0 dp_source2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .bus_readdatavalid_in(readmaster2_readdatavalid_in),
    .bus_readdatavalid_vm_in(readmaster2_readdatavalid_vm_in),
    .bus_readdata_in(readmaster2_readdata_in),
    .bus_wait_request_in(readmaster2_wait_request_in),
    .gen_valid_in(gen_sram_src_valid),
    .gen_vm_in(gen_sram_vm),
    .gen_fork_in(gen_sram_fork),
    .gen_data_flow_in(gen_sram_data_flow),
    .gen_src_stream_in(gen_sram_src_stream),
    .gen_dest_stream_in(gen_sram_dest_stream),
    .gen_stream_id_in(gen_sram_stream_id),
    .gen_src_vector_in(gen_sram_src_vector),
    .gen_dst_vector_in(gen_sram_dst_vector),
    .gen_src_scatter_in(gen_sram_src_scatter),
    .gen_dst_scatter_in(gen_sram_dst_scatter),
    .gen_src_start_in(gen_sram_src_start),
    .gen_src_end_in(gen_sram_src_end),
    .gen_dst_end_in(gen_sram_dst_end),
    .gen_src_eof_in(gen_sram_src_eof),
    .gen_src_addr_in(gen_sram_src_addr),
    .gen_src_addr_mode_in(gen_sram_src_addr_mode),
    .gen_dst_addr_in(gen_sram_dst_addr),
    .gen_dst_addr_mode_in(gen_sram_dst_addr_mode),
    .gen_bus_id_source_in(gen_sram_bus_id_source),
    .gen_data_type_source_in(gen_sram_data_type_source),
    .gen_data_model_source_in(gen_sram_data_model_source),
    .gen_bus_id_dest_in(gen_sram_bus_id_dest),
    .gen_busy_dest_in(gen_sram_busy_dest),
    .gen_data_type_dest_in(gen_sram_data_type_dest),
    .gen_data_model_dest_in(gen_sram_data_model_dest),
    .gen_src_burstlen_in(gen_sram_src_burstlen),
    .gen_dst_burstlen_in(gen_sram_dst_burstlen),
    .gen_thread_in(gen_sram_thread),
    .gen_mcast_in(gen_sram_mcast),
    .gen_src_data_in(gen_sram_data),
    .wr_full_in(n5707_o),
    .bus_addr_out(dp_source2_i_bus_addr_out),
    .bus_addr_mode_out(),
    .bus_cs_out(dp_source2_i_bus_cs_out),
    .bus_read_out(dp_source2_i_bus_read_out),
    .bus_read_vm_out(dp_source2_i_bus_read_vm_out),
    .bus_read_fork_out(dp_source2_i_bus_read_fork_out),
    .bus_read_data_flow_out(),
    .bus_read_stream_out(),
    .bus_read_stream_id_out(),
    .bus_read_vector_out(dp_source2_i_bus_read_vector_out),
    .bus_read_scatter_out(dp_source2_i_bus_read_scatter_out),
    .bus_read_start_out(),
    .bus_read_end_out(),
    .bus_burstlen_out(dp_source2_i_bus_burstlen_out),
    .bus_id_out(dp_source2_i_bus_id_out),
    .bus_data_type_out(),
    .bus_data_model_out(),
    .gen_waitreq_out(dp_source2_i_gen_waitreq_out),
    .wr_req_out(dp_source2_i_wr_req_out),
    .wr_req_pending_p0_out(dp_source2_i_wr_req_pending_p0_out),
    .wr_req_pending_p1_out(dp_source2_i_wr_req_pending_p1_out),
    .wr_data_flow_out(dp_source2_i_wr_data_flow_out),
    .wr_vector_out(dp_source2_i_wr_vector_out),
    .wr_stream_out(dp_source2_i_wr_stream_out),
    .wr_stream_id_out(dp_source2_i_wr_stream_id_out),
    .wr_scatter_out(dp_source2_i_wr_scatter_out),
    .wr_end_out(dp_source2_i_wr_end_out),
    .wr_addr_out(dp_source2_i_wr_addr_out),
    .wr_fork_out(dp_source2_i_wr_fork_out),
    .wr_addr_mode_out(dp_source2_i_wr_addr_mode_out),
    .wr_src_vm_out(dp_source2_i_wr_src_vm_out),
    .wr_datavalid_out(dp_source2_i_wr_datavalid_out),
    .wr_data_out(dp_source2_i_wr_data_out),
    .wr_readdatavalid_out(dp_source2_i_wr_readdatavalid_out),
    .wr_readdatavalid_vm_out(dp_source2_i_wr_readdatavalid_vm_out),
    .wr_readdata_out(dp_source2_i_wr_readdata_out),
    .wr_burstlen_out(dp_source2_i_wr_burstlen_out),
    .wr_bus_id_out(dp_source2_i_wr_bus_id_out),
    .wr_thread_out(dp_source2_i_wr_thread_out),
    .wr_data_type_out(dp_source2_i_wr_data_type_out),
    .wr_data_model_out(dp_source2_i_wr_data_model_out),
    .wr_mcast_out(dp_source2_i_wr_mcast_out));
  assign n5782_o = dp_source2_i_n5704[0];
  assign n5783_o = dp_source2_i_n5704[1];
  assign n5784_o = dp_source2_i_n5704[2];
  assign n5786_o = dp_source2_i_n5705[0];
  assign n5787_o = dp_source2_i_n5705[1];
  assign n5788_o = dp_source2_i_n5705[2];
  assign n5790_o = dp_source2_i_n5706[0];
  assign n5791_o = dp_source2_i_n5706[1];
  assign n5792_o = dp_source2_i_n5706[2];
  assign n5794_o = dp_source2_i_n5708[1:0];
  assign n5795_o = dp_source2_i_n5708[3:2];
  assign n5796_o = dp_source2_i_n5708[5:4];
  assign n5798_o = dp_source2_i_n5709[2:0];
  assign n5799_o = dp_source2_i_n5709[5:3];
  assign n5800_o = dp_source2_i_n5709[8:6];
  assign n5802_o = dp_source2_i_n5710[0];
  assign n5806_o = dp_source2_i_n5711[1:0];
  assign n5810_o = dp_source2_i_n5712[1:0];
  assign n5811_o = dp_source2_i_n5712[3:2];
  assign n5812_o = dp_source2_i_n5712[5:4];
  assign n5814_o = dp_source2_i_n5713[3:0];
  assign n5815_o = dp_source2_i_n5713[7:4];
  assign n5816_o = dp_source2_i_n5713[11:8];
  /* ../../HW/src/dp/dp.vhd:910:27  */
  assign dp_source3_i0_n5832 = dp_source3_i0_bus_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:911:25  */
  assign dp_source3_i0_n5834 = dp_source3_i0_bus_cs_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:912:27  */
  assign dp_source3_i0_n5835 = dp_source3_i0_bus_read_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:913:30  */
  assign dp_source3_i0_n5836 = dp_source3_i0_bus_read_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:918:34  */
  assign dp_source3_i0_n5841 = dp_source3_i0_bus_read_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:919:35  */
  assign dp_source3_i0_n5842 = dp_source3_i0_bus_read_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:920:33  */
  assign dp_source3_i0_n5843 = dp_source3_i0_bus_read_start_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:921:31  */
  assign dp_source3_i0_n5844 = dp_source3_i0_bus_read_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:926:31  */
  assign dp_source3_i0_n5845 = dp_source3_i0_bus_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:927:25  */
  assign dp_source3_i0_n5846 = dp_source3_i0_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:931:30  */
  assign dp_source3_i0_n5849 = dp_source3_i0_gen_waitreq_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:964:29  */
  assign dp_source3_i0_n5850 = dp_source3_i0_wr_req_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:968:40  */
  assign dp_source3_i0_n5851 = dp_source3_i0_wr_req_pending_p0_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:972:40  */
  assign dp_source3_i0_n5852 = dp_source3_i0_wr_req_pending_p1_out; // (signal)
  assign n5853_o = {wr_ddr_full, wr_sram_full, wr_full};
  /* ../../HW/src/dp/dp.vhd:980:34  */
  assign dp_source3_i0_n5854 = dp_source3_i0_wr_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:992:31  */
  assign dp_source3_i0_n5855 = dp_source3_i0_wr_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:984:31  */
  assign dp_source3_i0_n5856 = dp_source3_i0_wr_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:988:34  */
  assign dp_source3_i0_n5857 = dp_source3_i0_wr_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:996:32  */
  assign dp_source3_i0_n5858 = dp_source3_i0_wr_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1000:28  */
  assign dp_source3_i0_n5859 = dp_source3_i0_wr_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1004:27  */
  assign dp_source3_i0_n5860 = dp_source3_i0_wr_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1006:27  */
  assign dp_source3_i0_n5861 = dp_source3_i0_wr_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1010:30  */
  assign dp_source3_i0_n5862 = dp_source3_i0_wr_src_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1008:31  */
  assign dp_source3_i0_n5863 = dp_source3_i0_wr_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1012:33  */
  assign dp_source3_i0_n5864 = dp_source3_i0_wr_datavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1014:27  */
  assign dp_source3_i0_n5865 = dp_source3_i0_wr_data_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1016:37  */
  assign dp_source3_i0_n5866 = dp_source3_i0_wr_readdatavalid_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1018:40  */
  assign dp_source3_i0_n5867 = dp_source3_i0_wr_readdatavalid_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1020:32  */
  assign dp_source3_i0_n5868 = dp_source3_i0_wr_readdata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1022:31  */
  assign dp_source3_i0_n5869 = dp_source3_i0_wr_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1024:29  */
  assign dp_source3_i0_n5870 = dp_source3_i0_wr_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1026:28  */
  assign dp_source3_i0_n5871 = dp_source3_i0_wr_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1028:31  */
  assign dp_source3_i0_n5872 = dp_source3_i0_wr_data_type_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1030:32  */
  assign dp_source3_i0_n5873 = dp_source3_i0_wr_data_model_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1032:27  */
  assign dp_source3_i0_n5874 = dp_source3_i0_wr_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:897:1  */
  dp_source_2_3_1_32_1_0 dp_source3_i0 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .bus_readdatavalid_in(readmaster3_readdatavalid_in),
    .bus_readdatavalid_vm_in(readmaster3_readdatavalid_vm_in),
    .bus_readdata_in(readmaster3_readdata_in),
    .bus_wait_request_in(readmaster3_wait_request_in),
    .gen_valid_in(gen_ddr_src_valid),
    .gen_vm_in(gen_ddr_vm),
    .gen_fork_in(gen_ddr_fork),
    .gen_data_flow_in(gen_ddr_data_flow),
    .gen_src_stream_in(gen_ddr_src_stream),
    .gen_dest_stream_in(gen_ddr_dest_stream),
    .gen_stream_id_in(gen_ddr_stream_id),
    .gen_src_vector_in(gen_ddr_src_vector),
    .gen_dst_vector_in(gen_ddr_dst_vector),
    .gen_src_scatter_in(gen_ddr_src_scatter),
    .gen_dst_scatter_in(gen_ddr_dst_scatter),
    .gen_src_start_in(gen_ddr_src_start),
    .gen_src_end_in(gen_ddr_src_end),
    .gen_dst_end_in(gen_ddr_dst_end),
    .gen_src_eof_in(gen_ddr_src_eof),
    .gen_src_addr_in(gen_ddr_src_addr),
    .gen_src_addr_mode_in(gen_ddr_src_addr_mode),
    .gen_dst_addr_in(gen_ddr_dst_addr),
    .gen_dst_addr_mode_in(gen_ddr_dst_addr_mode),
    .gen_bus_id_source_in(gen_ddr_bus_id_source),
    .gen_data_type_source_in(gen_ddr_data_type_source),
    .gen_data_model_source_in(gen_ddr_data_model_source),
    .gen_bus_id_dest_in(gen_ddr_bus_id_dest),
    .gen_busy_dest_in(gen_ddr_busy_dest),
    .gen_data_type_dest_in(gen_ddr_data_type_dest),
    .gen_data_model_dest_in(gen_ddr_data_model_dest),
    .gen_src_burstlen_in(gen_ddr_src_burstlen),
    .gen_dst_burstlen_in(gen_ddr_dst_burstlen),
    .gen_thread_in(gen_ddr_thread),
    .gen_mcast_in(gen_ddr_mcast),
    .gen_src_data_in(gen_ddr_data),
    .wr_full_in(n5853_o),
    .bus_addr_out(dp_source3_i0_bus_addr_out),
    .bus_addr_mode_out(),
    .bus_cs_out(dp_source3_i0_bus_cs_out),
    .bus_read_out(dp_source3_i0_bus_read_out),
    .bus_read_vm_out(dp_source3_i0_bus_read_vm_out),
    .bus_read_fork_out(),
    .bus_read_data_flow_out(),
    .bus_read_stream_out(),
    .bus_read_stream_id_out(),
    .bus_read_vector_out(dp_source3_i0_bus_read_vector_out),
    .bus_read_scatter_out(dp_source3_i0_bus_read_scatter_out),
    .bus_read_start_out(dp_source3_i0_bus_read_start_out),
    .bus_read_end_out(dp_source3_i0_bus_read_end_out),
    .bus_burstlen_out(dp_source3_i0_bus_burstlen_out),
    .bus_id_out(dp_source3_i0_bus_id_out),
    .bus_data_type_out(),
    .bus_data_model_out(),
    .gen_waitreq_out(dp_source3_i0_gen_waitreq_out),
    .wr_req_out(dp_source3_i0_wr_req_out),
    .wr_req_pending_p0_out(dp_source3_i0_wr_req_pending_p0_out),
    .wr_req_pending_p1_out(dp_source3_i0_wr_req_pending_p1_out),
    .wr_data_flow_out(dp_source3_i0_wr_data_flow_out),
    .wr_vector_out(dp_source3_i0_wr_vector_out),
    .wr_stream_out(dp_source3_i0_wr_stream_out),
    .wr_stream_id_out(dp_source3_i0_wr_stream_id_out),
    .wr_scatter_out(dp_source3_i0_wr_scatter_out),
    .wr_end_out(dp_source3_i0_wr_end_out),
    .wr_addr_out(dp_source3_i0_wr_addr_out),
    .wr_fork_out(dp_source3_i0_wr_fork_out),
    .wr_addr_mode_out(dp_source3_i0_wr_addr_mode_out),
    .wr_src_vm_out(dp_source3_i0_wr_src_vm_out),
    .wr_datavalid_out(dp_source3_i0_wr_datavalid_out),
    .wr_data_out(dp_source3_i0_wr_data_out),
    .wr_readdatavalid_out(dp_source3_i0_wr_readdatavalid_out),
    .wr_readdatavalid_vm_out(dp_source3_i0_wr_readdatavalid_vm_out),
    .wr_readdata_out(dp_source3_i0_wr_readdata_out),
    .wr_burstlen_out(dp_source3_i0_wr_burstlen_out),
    .wr_bus_id_out(dp_source3_i0_wr_bus_id_out),
    .wr_thread_out(dp_source3_i0_wr_thread_out),
    .wr_data_type_out(dp_source3_i0_wr_data_type_out),
    .wr_data_model_out(dp_source3_i0_wr_data_model_out),
    .wr_mcast_out(dp_source3_i0_wr_mcast_out));
  assign n5929_o = dp_source3_i0_n5850[0];
  assign n5930_o = dp_source3_i0_n5850[1];
  assign n5931_o = dp_source3_i0_n5850[2];
  assign n5933_o = dp_source3_i0_n5851[0];
  assign n5934_o = dp_source3_i0_n5851[1];
  assign n5935_o = dp_source3_i0_n5851[2];
  assign n5937_o = dp_source3_i0_n5852[0];
  assign n5938_o = dp_source3_i0_n5852[1];
  assign n5939_o = dp_source3_i0_n5852[2];
  assign n5941_o = dp_source3_i0_n5854[1:0];
  assign n5942_o = dp_source3_i0_n5854[3:2];
  assign n5943_o = dp_source3_i0_n5854[5:4];
  assign n5945_o = dp_source3_i0_n5855[2:0];
  assign n5946_o = dp_source3_i0_n5855[5:3];
  assign n5947_o = dp_source3_i0_n5855[8:6];
  assign n5949_o = dp_source3_i0_n5856[0];
  assign n5953_o = dp_source3_i0_n5857[1:0];
  assign n5957_o = dp_source3_i0_n5858[1:0];
  assign n5958_o = dp_source3_i0_n5858[3:2];
  assign n5959_o = dp_source3_i0_n5858[5:4];
  assign n5961_o = dp_source3_i0_n5859[3:0];
  assign n5962_o = dp_source3_i0_n5859[7:4];
  assign n5963_o = dp_source3_i0_n5859[11:8];
  /* ../../HW/src/dp/dp.vhd:1052:27  */
  assign dp_sink1_i_n5979 = dp_sink1_i_bus_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1053:27  */
  assign dp_sink1_i_n5980 = dp_sink1_i_bus_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1054:32  */
  assign dp_sink1_i_n5981 = dp_sink1_i_bus_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1055:25  */
  assign dp_sink1_i_n5982 = dp_sink1_i_bus_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1056:32  */
  assign dp_sink1_i_n5983 = dp_sink1_i_bus_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1057:29  */
  assign dp_sink1_i_n5984 = dp_sink1_i_bus_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1058:29  */
  assign dp_sink1_i_n5985 = dp_sink1_i_bus_stream_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1059:32  */
  assign dp_sink1_i_n5986 = dp_sink1_i_bus_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1060:30  */
  assign dp_sink1_i_n5987 = dp_sink1_i_bus_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1062:28  */
  assign dp_sink1_i_n5989 = dp_sink1_i_bus_mcast_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1063:25  */
  assign dp_sink1_i_n5990 = dp_sink1_i_bus_cs_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1064:28  */
  assign dp_sink1_i_n5991 = dp_sink1_i_bus_write_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1065:32  */
  assign dp_sink1_i_n5992 = dp_sink1_i_bus_writedata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1067:31  */
  assign dp_sink1_i_n5993 = dp_sink1_i_bus_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1070:25  */
  assign dp_sink1_i_n5996 = dp_sink1_i_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1071:32  */
  assign dp_sink1_i_n5997 = dp_sink1_i_bus_data_type_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1072:33  */
  assign dp_sink1_i_n5998 = dp_sink1_i_bus_data_model_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1073:29  */
  assign dp_sink1_i_n5999 = dp_sink1_i_bus_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1075:34  */
  assign dp_sink1_i_n6000 = dp_sink1_i_wr_maxburstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1076:27  */
  assign dp_sink1_i_n6001 = dp_sink1_i_wr_full_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1102:34  */
  assign dp_sink1_i_n6002 = dp_sink1_i_read_pending_p0_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1103:34  */
  assign dp_sink1_i_n6003 = dp_sink1_i_read_pending_p1_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1040:1  */
  dp_sink_3_32_1_9_6a0e3f59309a30c5143aeb870000c064ad45653d dp_sink1_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .bus_wait_request_in(writemaster1_wait_request_in),
    .wr_req_in(wr_req),
    .wr_req_pending_p0_in(wr_req_p0_pending),
    .wr_req_pending_p1_in(wr_req_p1_pending),
    .wr_data_flow_in(wr_data_flow),
    .wr_vector_in(wr_vector),
    .wr_stream_in(wr_stream),
    .wr_stream_id_in(wr_stream_id),
    .wr_scatter_in(wr_scatter),
    .wr_end_in(wr_end),
    .wr_addr_in(wr_addr),
    .wr_fork_in(wr_fork),
    .wr_addr_mode_in(wr_addr_mode),
    .wr_src_vm_in(wr_src_vm),
    .wr_datavalid_in(wr_datavalid),
    .wr_data_in(wr_data),
    .wr_readdatavalid_in(wr_readdatavalid),
    .wr_readdatavalid_vm_in(wr_readdatavalid_vm),
    .wr_readdata_in(wr_readdata),
    .wr_burstlen_in(wr_burstlen),
    .wr_bus_id_in(wr_bus_id),
    .wr_thread_in(wr_thread),
    .wr_data_type_in(wr_data_type),
    .wr_data_model_in(wr_data_model),
    .wr_mcast_in(wr_mcast),
    .bus_addr_out(dp_sink1_i_bus_addr_out),
    .bus_fork_out(dp_sink1_i_bus_fork_out),
    .bus_addr_mode_out(dp_sink1_i_bus_addr_mode_out),
    .bus_vm_out(dp_sink1_i_bus_vm_out),
    .bus_data_flow_out(dp_sink1_i_bus_data_flow_out),
    .bus_vector_out(dp_sink1_i_bus_vector_out),
    .bus_stream_out(dp_sink1_i_bus_stream_out),
    .bus_stream_id_out(dp_sink1_i_bus_stream_id_out),
    .bus_scatter_out(dp_sink1_i_bus_scatter_out),
    .bus_end_out(),
    .bus_mcast_out(dp_sink1_i_bus_mcast_out),
    .bus_cs_out(dp_sink1_i_bus_cs_out),
    .bus_write_out(dp_sink1_i_bus_write_out),
    .bus_writedata_out(dp_sink1_i_bus_writedata_out),
    .bus_burstlen_out(dp_sink1_i_bus_burstlen_out),
    .bus_burstlen2_out(),
    .bus_burstlen3_out(),
    .bus_id_out(dp_sink1_i_bus_id_out),
    .bus_data_type_out(dp_sink1_i_bus_data_type_out),
    .bus_data_model_out(dp_sink1_i_bus_data_model_out),
    .bus_thread_out(dp_sink1_i_bus_thread_out),
    .wr_maxburstlen_out(dp_sink1_i_wr_maxburstlen_out),
    .wr_full_out(dp_sink1_i_wr_full_out),
    .read_pending_p0_out(dp_sink1_i_read_pending_p0_out),
    .read_pending_p1_out(dp_sink1_i_read_pending_p1_out));
  /* ../../HW/src/dp/dp.vhd:1122:27  */
  assign dp_sink2_i_n6051 = dp_sink2_i_bus_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1123:27  */
  assign dp_sink2_i_n6052 = dp_sink2_i_bus_fork_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1125:25  */
  assign dp_sink2_i_n6054 = dp_sink2_i_bus_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1127:29  */
  assign dp_sink2_i_n6056 = dp_sink2_i_bus_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1130:30  */
  assign dp_sink2_i_n6059 = dp_sink2_i_bus_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1133:25  */
  assign dp_sink2_i_n6062 = dp_sink2_i_bus_cs_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1134:28  */
  assign dp_sink2_i_n6063 = dp_sink2_i_bus_write_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1135:32  */
  assign dp_sink2_i_n6064 = dp_sink2_i_bus_writedata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1137:31  */
  assign dp_sink2_i_n6065 = dp_sink2_i_bus_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1140:25  */
  assign dp_sink2_i_n6068 = dp_sink2_i_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1143:29  */
  assign dp_sink2_i_n6071 = dp_sink2_i_bus_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1145:34  */
  assign dp_sink2_i_n6072 = dp_sink2_i_wr_maxburstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1146:27  */
  assign dp_sink2_i_n6073 = dp_sink2_i_wr_full_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1171:34  */
  assign dp_sink2_i_n6076 = dp_sink2_i_read_pending_p0_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1172:34  */
  assign dp_sink2_i_n6077 = dp_sink2_i_read_pending_p1_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1110:1  */
  dp_sink_3_32_1_9_6a0e3f59309a30c5143aeb870000c064ad45653d dp_sink2_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .bus_wait_request_in(writemaster2_wait_request_in),
    .wr_req_in(wr_sram_req),
    .wr_req_pending_p0_in(wr_sram_req_p0_pending),
    .wr_req_pending_p1_in(wr_sram_req_p1_pending),
    .wr_data_flow_in(wr_sram_data_flow),
    .wr_vector_in(wr_sram_vector),
    .wr_stream_in(n6074_o),
    .wr_stream_id_in(n6075_o),
    .wr_scatter_in(wr_sram_scatter),
    .wr_end_in(wr_sram_end),
    .wr_addr_in(wr_addr),
    .wr_fork_in(wr_fork),
    .wr_addr_mode_in(wr_addr_mode),
    .wr_src_vm_in(wr_src_vm),
    .wr_datavalid_in(wr_datavalid),
    .wr_data_in(wr_data),
    .wr_readdatavalid_in(wr_readdatavalid),
    .wr_readdatavalid_vm_in(wr_readdatavalid_vm),
    .wr_readdata_in(wr_readdata),
    .wr_burstlen_in(wr_burstlen),
    .wr_bus_id_in(wr_bus_id),
    .wr_thread_in(wr_thread),
    .wr_data_type_in(wr_data_type),
    .wr_data_model_in(wr_data_model),
    .wr_mcast_in(wr_mcast),
    .bus_addr_out(dp_sink2_i_bus_addr_out),
    .bus_fork_out(dp_sink2_i_bus_fork_out),
    .bus_addr_mode_out(),
    .bus_vm_out(dp_sink2_i_bus_vm_out),
    .bus_data_flow_out(),
    .bus_vector_out(dp_sink2_i_bus_vector_out),
    .bus_stream_out(),
    .bus_stream_id_out(),
    .bus_scatter_out(dp_sink2_i_bus_scatter_out),
    .bus_end_out(),
    .bus_mcast_out(),
    .bus_cs_out(dp_sink2_i_bus_cs_out),
    .bus_write_out(dp_sink2_i_bus_write_out),
    .bus_writedata_out(dp_sink2_i_bus_writedata_out),
    .bus_burstlen_out(dp_sink2_i_bus_burstlen_out),
    .bus_burstlen2_out(),
    .bus_burstlen3_out(),
    .bus_id_out(dp_sink2_i_bus_id_out),
    .bus_data_type_out(),
    .bus_data_model_out(),
    .bus_thread_out(dp_sink2_i_bus_thread_out),
    .wr_maxburstlen_out(dp_sink2_i_wr_maxburstlen_out),
    .wr_full_out(dp_sink2_i_wr_full_out),
    .read_pending_p0_out(dp_sink2_i_read_pending_p0_out),
    .read_pending_p1_out(dp_sink2_i_read_pending_p1_out));
  /* ../../HW/src/dp/dp.vhd:1191:27  */
  assign dp_sink3_i_n6118 = dp_sink3_i_bus_addr_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1194:25  */
  assign dp_sink3_i_n6121 = dp_sink3_i_bus_vm_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1196:29  */
  assign dp_sink3_i_n6123 = dp_sink3_i_bus_vector_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1199:30  */
  assign dp_sink3_i_n6126 = dp_sink3_i_bus_scatter_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1200:26  */
  assign dp_sink3_i_n6127 = dp_sink3_i_bus_end_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1202:25  */
  assign dp_sink3_i_n6129 = dp_sink3_i_bus_cs_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1203:28  */
  assign dp_sink3_i_n6130 = dp_sink3_i_bus_write_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1204:32  */
  assign dp_sink3_i_n6131 = dp_sink3_i_bus_writedata_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1206:31  */
  assign dp_sink3_i_n6132 = dp_sink3_i_bus_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1207:32  */
  assign dp_sink3_i_n6133 = dp_sink3_i_bus_burstlen2_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1208:32  */
  assign dp_sink3_i_n6134 = dp_sink3_i_bus_burstlen3_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1209:25  */
  assign dp_sink3_i_n6135 = dp_sink3_i_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1212:29  */
  assign dp_sink3_i_n6138 = dp_sink3_i_bus_thread_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1214:34  */
  assign dp_sink3_i_n6139 = dp_sink3_i_wr_maxburstlen_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1215:27  */
  assign dp_sink3_i_n6140 = dp_sink3_i_wr_full_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1240:34  */
  assign dp_sink3_i_n6143 = dp_sink3_i_read_pending_p0_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1241:34  */
  assign dp_sink3_i_n6144 = dp_sink3_i_read_pending_p1_out; // (signal)
  /* ../../HW/src/dp/dp.vhd:1179:1  */
  dp_sink_3_32_1_9_40623dc9948b5e96ae4a8c3b66bafc8116c42db3 dp_sink3_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .bus_wait_request_in(writemaster3_wait_request_in),
    .wr_req_in(wr_ddr_req),
    .wr_req_pending_p0_in(wr_ddr_req_p0_pending),
    .wr_req_pending_p1_in(wr_ddr_req_p1_pending),
    .wr_data_flow_in(wr_ddr_data_flow),
    .wr_vector_in(wr_ddr_vector),
    .wr_stream_in(n6141_o),
    .wr_stream_id_in(n6142_o),
    .wr_scatter_in(wr_ddr_scatter),
    .wr_end_in(wr_ddr_end),
    .wr_addr_in(wr_addr),
    .wr_fork_in(wr_fork),
    .wr_addr_mode_in(wr_addr_mode),
    .wr_src_vm_in(wr_src_vm),
    .wr_datavalid_in(wr_datavalid),
    .wr_data_in(wr_data),
    .wr_readdatavalid_in(wr_readdatavalid),
    .wr_readdatavalid_vm_in(wr_readdatavalid_vm),
    .wr_readdata_in(wr_readdata),
    .wr_burstlen_in(wr_burstlen),
    .wr_bus_id_in(wr_bus_id),
    .wr_thread_in(wr_thread),
    .wr_data_type_in(wr_data_type),
    .wr_data_model_in(wr_data_model),
    .wr_mcast_in(wr_mcast),
    .bus_addr_out(dp_sink3_i_bus_addr_out),
    .bus_fork_out(),
    .bus_addr_mode_out(),
    .bus_vm_out(dp_sink3_i_bus_vm_out),
    .bus_data_flow_out(),
    .bus_vector_out(dp_sink3_i_bus_vector_out),
    .bus_stream_out(),
    .bus_stream_id_out(),
    .bus_scatter_out(dp_sink3_i_bus_scatter_out),
    .bus_end_out(dp_sink3_i_bus_end_out),
    .bus_mcast_out(),
    .bus_cs_out(dp_sink3_i_bus_cs_out),
    .bus_write_out(dp_sink3_i_bus_write_out),
    .bus_writedata_out(dp_sink3_i_bus_writedata_out),
    .bus_burstlen_out(dp_sink3_i_bus_burstlen_out),
    .bus_burstlen2_out(dp_sink3_i_bus_burstlen2_out),
    .bus_burstlen3_out(dp_sink3_i_bus_burstlen3_out),
    .bus_id_out(dp_sink3_i_bus_id_out),
    .bus_data_type_out(),
    .bus_data_model_out(),
    .bus_thread_out(dp_sink3_i_bus_thread_out),
    .wr_maxburstlen_out(dp_sink3_i_wr_maxburstlen_out),
    .wr_full_out(dp_sink3_i_wr_full_out),
    .read_pending_p0_out(dp_sink3_i_read_pending_p0_out),
    .read_pending_p1_out(dp_sink3_i_read_pending_p1_out));
  assign n6187_o = {dp_source3_i0_n5864, dp_source2_i_n5718, dp_source1_i_n5566};
  assign n6188_o = {dp_source3_i0_n5860, dp_source2_i_n5714, dp_source1_i_n5562};
  assign n6189_o = {dp_source3_i0_n5861, dp_source2_i_n5715, dp_source1_i_n5563};
  assign n6190_o = {dp_source3_i0_n5863, dp_source2_i_n5717, dp_source1_i_n5565};
  assign n6191_o = {dp_source3_i0_n5862, dp_source2_i_n5716, dp_source1_i_n5564};
  assign n6192_o = {dp_source3_i0_n5865, dp_source2_i_n5719, dp_source1_i_n5567};
  assign n6193_o = {dp_source3_i0_n5868, dp_source2_i_n5722, dp_source1_i_n5570};
  assign n6194_o = {dp_source3_i0_n5866, dp_source2_i_n5720, dp_source1_i_n5568};
  assign n6195_o = {dp_source3_i0_n5867, dp_source2_i_n5721, dp_source1_i_n5569};
  assign n6196_o = {dp_source3_i0_n5869, dp_source2_i_n5723, dp_source1_i_n5571};
  assign n6197_o = {dp_source3_i0_n5870, dp_source2_i_n5724, dp_source1_i_n5572};
  assign n6198_o = {dp_source3_i0_n5871, dp_source2_i_n5725, dp_source1_i_n5573};
  assign n6199_o = {dp_source3_i0_n5872, dp_source2_i_n5726, dp_source1_i_n5574};
  assign n6200_o = {dp_source3_i0_n5873, dp_source2_i_n5727, dp_source1_i_n5575};
  assign n6201_o = {dp_source3_i0_n5874, dp_source2_i_n5728, dp_source1_i_n5576};
  assign n6202_o = {dp_source3_i0_n5849, dp_source2_i_n5703, dp_source1_i_n5551};
  assign n6203_o = {n5929_o, n5782_o, n5636_o};
  assign n6204_o = {n5933_o, n5786_o, n5640_o};
  assign n6205_o = {n5937_o, n5790_o, n5644_o};
  assign n6206_o = {n5930_o, n5783_o, n5637_o};
  assign n6207_o = {n5934_o, n5787_o, n5641_o};
  assign n6208_o = {n5938_o, n5791_o, n5645_o};
  assign n6209_o = {n5931_o, n5784_o, n5638_o};
  assign n6210_o = {n5935_o, n5788_o, n5642_o};
  assign n6211_o = {n5939_o, n5792_o, n5646_o};
  assign n6226_o = {wr_ddr_full, wr_sram_full, wr_full};
  assign n6227_o = {dp_sink3_i_n6139, dp_sink2_i_n6072, dp_sink1_i_n6000};
  assign n6228_o = {n5945_o, n5798_o, n5652_o};
  assign n6229_o = {n5946_o, n5799_o, n5653_o};
  assign n6230_o = {n5947_o, n5800_o, n5654_o};
  assign n6231_o = {n5957_o, n5810_o, n5664_o};
  assign n6232_o = {n5958_o, n5811_o, n5665_o};
  assign n6233_o = {n5959_o, n5812_o, n5666_o};
  assign n6234_o = {n5961_o, n5814_o, n5668_o};
  assign n6235_o = {n5962_o, n5815_o, n5669_o};
  assign n6236_o = {n5963_o, n5816_o, n5670_o};
  assign n6237_o = {n5941_o, n5794_o, n5648_o};
  assign n6238_o = {n5942_o, n5795_o, n5649_o};
  assign n6239_o = {n5943_o, n5796_o, n5650_o};
  assign n6240_o = {n5949_o, n5802_o, n5656_o};
  assign n6243_o = {n5953_o, n5806_o, n5660_o};
endmodule

module scfifo_35_6_53_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [34:0] data_in,
   input  write_in,
   input  read_in,
   output [34:0] q_out,
   output [5:0] ravail_out,
   output [5:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [34:0] q;
  wire [5:0] address_a;
  wire [5:0] address_b;
  wire [5:0] waddr_r;
  wire [5:0] waddr_rr;
  wire [5:0] raddr_r;
  wire [5:0] raddr;
  wire [5:0] ravail;
  wire [5:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [34:0] ram_i_n4989;
  wire [34:0] ram_i_q_b;
  wire [5:0] n4992_o;
  wire [5:0] n4993_o;
  wire n4994_o;
  wire n4997_o;
  wire n4998_o;
  wire [5:0] n5001_o;
  wire [5:0] n5002_o;
  wire n5005_o;
  wire [5:0] n5008_o;
  wire [5:0] n5010_o;
  wire n5011_o;
  wire n5014_o;
  wire [5:0] n5016_o;
  wire n5017_o;
  wire n5020_o;
  wire n5022_o;
  wire n5024_o;
  wire n5027_o;
  wire [5:0] n5049_o;
  reg [5:0] n5050_q;
  reg [5:0] n5051_q;
  reg [5:0] n5052_q;
  reg n5054_q;
  reg n5055_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n4994_o;
  assign full_out = full_r;
  assign almost_full_out = n4998_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n4989; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n5050_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n5051_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n5052_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n5002_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n4992_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n4993_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n5054_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n5055_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n4989 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_64_64_6_6_35_35 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n4992_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n4993_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n4994_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n4997_o = $unsigned(wused) >= $unsigned(6'b110101);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n4998_o = n4997_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n5001_o = raddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n5002_o = read_in ? n5001_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n5005_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n5008_o = waddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n5010_o = waddr_r + 6'b000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n5011_o = n5010_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n5014_o = n5011_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n5016_o = waddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n5017_o = n5016_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n5020_o = n5017_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n5022_o = write_in ? n5014_o : n5020_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n5024_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n5027_o = n5024_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n5049_o = write_in ? n5008_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n5005_o)
    if (n5005_o)
      n5050_q <= 6'b000000;
    else
      n5050_q <= n5049_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n5005_o)
    if (n5005_o)
      n5051_q <= 6'b000000;
    else
      n5051_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n5005_o)
    if (n5005_o)
      n5052_q <= 6'b000000;
    else
      n5052_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n5005_o)
    if (n5005_o)
      n5054_q <= 1'b0;
    else
      n5054_q <= n5027_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n5005_o)
    if (n5005_o)
      n5055_q <= 1'b0;
    else
      n5055_q <= n5022_o;
endmodule

module scfifo_37_4_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [36:0] data_in,
   input  write_in,
   input  read_in,
   output [36:0] q_out,
   output [3:0] ravail_out,
   output [3:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [36:0] q;
  wire [3:0] address_a;
  wire [3:0] address_b;
  wire [3:0] waddr_r;
  wire [3:0] waddr_rr;
  wire [3:0] raddr_r;
  wire [3:0] raddr;
  wire [3:0] ravail;
  wire [3:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [36:0] ram_i_n4916;
  wire [36:0] ram_i_q_b;
  wire [3:0] n4919_o;
  wire [3:0] n4920_o;
  wire n4921_o;
  wire n4924_o;
  wire n4925_o;
  wire [3:0] n4928_o;
  wire [3:0] n4929_o;
  wire n4932_o;
  wire [3:0] n4935_o;
  wire [3:0] n4937_o;
  wire n4938_o;
  wire n4941_o;
  wire [3:0] n4943_o;
  wire n4944_o;
  wire n4947_o;
  wire n4949_o;
  wire n4951_o;
  wire n4954_o;
  wire [3:0] n4976_o;
  reg [3:0] n4977_q;
  reg [3:0] n4978_q;
  reg [3:0] n4979_q;
  reg n4981_q;
  reg n4982_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n4921_o;
  assign full_out = full_r;
  assign almost_full_out = n4925_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n4916; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n4977_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n4978_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n4979_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n4929_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n4919_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n4920_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n4981_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n4982_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n4916 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_16_16_4_4_37_37 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n4919_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n4920_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n4921_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n4924_o = $unsigned(wused) >= $unsigned(4'b0001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n4925_o = n4924_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n4928_o = raddr_r + 4'b0001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n4929_o = read_in ? n4928_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n4932_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n4935_o = waddr_r + 4'b0001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n4937_o = waddr_r + 4'b0010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n4938_o = n4937_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n4941_o = n4938_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n4943_o = waddr_r + 4'b0001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n4944_o = n4943_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n4947_o = n4944_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n4949_o = write_in ? n4941_o : n4947_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n4951_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n4954_o = n4951_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n4976_o = write_in ? n4935_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4932_o)
    if (n4932_o)
      n4977_q <= 4'b0000;
    else
      n4977_q <= n4976_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4932_o)
    if (n4932_o)
      n4978_q <= 4'b0000;
    else
      n4978_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4932_o)
    if (n4932_o)
      n4979_q <= 4'b0000;
    else
      n4979_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4932_o)
    if (n4932_o)
      n4981_q <= 1'b0;
    else
      n4981_q <= n4954_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4932_o)
    if (n4932_o)
      n4982_q <= 1'b0;
    else
      n4982_q <= n4949_o;
endmodule

module scfifo_64_9_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [63:0] data_in,
   input  write_in,
   input  read_in,
   output [63:0] q_out,
   output [8:0] ravail_out,
   output [8:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [63:0] q;
  wire [8:0] address_a;
  wire [8:0] address_b;
  wire [8:0] waddr_r;
  wire [8:0] waddr_rr;
  wire [8:0] raddr_r;
  wire [8:0] raddr;
  wire [8:0] ravail;
  wire [8:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [63:0] ram_i_n4843;
  wire [63:0] ram_i_q_b;
  wire [8:0] n4846_o;
  wire [8:0] n4847_o;
  wire n4848_o;
  wire n4851_o;
  wire n4852_o;
  wire [8:0] n4855_o;
  wire [8:0] n4856_o;
  wire n4859_o;
  wire [8:0] n4862_o;
  wire [8:0] n4864_o;
  wire n4865_o;
  wire n4868_o;
  wire [8:0] n4870_o;
  wire n4871_o;
  wire n4874_o;
  wire n4876_o;
  wire n4878_o;
  wire n4881_o;
  wire [8:0] n4903_o;
  reg [8:0] n4904_q;
  reg [8:0] n4905_q;
  reg [8:0] n4906_q;
  reg n4908_q;
  reg n4909_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n4848_o;
  assign full_out = full_r;
  assign almost_full_out = n4852_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n4843; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n4904_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n4905_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n4906_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n4856_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n4846_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n4847_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n4908_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n4909_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n4843 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_512_512_9_9_64_64 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n4846_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n4847_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n4848_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n4851_o = $unsigned(wused) >= $unsigned(9'b000000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n4852_o = n4851_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n4855_o = raddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n4856_o = read_in ? n4855_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n4859_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n4862_o = waddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n4864_o = waddr_r + 9'b000000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n4865_o = n4864_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n4868_o = n4865_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n4870_o = waddr_r + 9'b000000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n4871_o = n4870_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n4874_o = n4871_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n4876_o = write_in ? n4868_o : n4874_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n4878_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n4881_o = n4878_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n4903_o = write_in ? n4862_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4859_o)
    if (n4859_o)
      n4904_q <= 9'b000000000;
    else
      n4904_q <= n4903_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4859_o)
    if (n4859_o)
      n4905_q <= 9'b000000000;
    else
      n4905_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4859_o)
    if (n4859_o)
      n4906_q <= 9'b000000000;
    else
      n4906_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4859_o)
    if (n4859_o)
      n4908_q <= 1'b0;
    else
      n4908_q <= n4881_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4859_o)
    if (n4859_o)
      n4909_q <= 1'b0;
    else
      n4909_q <= n4876_o;
endmodule

module sram_14
  (input  clock_in,
   input  reset_in,
   input  [13:0] dp_rd_addr_in,
   input  [13:0] dp_wr_addr_in,
   input  dp_write_in,
   input  [2:0] dp_write_vector_in,
   input  dp_read_in,
   input  [2:0] dp_read_vector_in,
   input  dp_read_gen_valid_in,
   input  [63:0] dp_writedata_in,
   output dp_readdatavalid_out,
   output [63:0] dp_readdata_out);
  wire [63:0] q;
  wire [63:0] q_r;
  wire rden_r;
  wire rden_rr;
  wire rden_rrr;
  wire [2:0] rd_vector_r;
  wire [2:0] rd_vector_rr;
  wire [2:0] rd_vector_rrr;
  wire valid;
  wire [10:0] dp_wr_addr;
  wire [13:0] rd_addr_r;
  wire [13:0] rd_addr_rr;
  wire [13:0] rd_addr_rrr;
  wire [7:0] byteena;
  wire [63:0] dp_writedata;
  wire [10:0] wr_addr_r;
  wire [7:0] byteena_r;
  wire [63:0] writedata_r;
  wire wren_r;
  wire [63:0] dp_readdata_r;
  wire dp_readdatavalid;
  wire dp_readdatavalid_r;
  wire n4519_o;
  wire delay_i1_n4522;
  localparam n4523_o = 1'b1;
  wire delay_i1_out_out;
  wire [10:0] n4526_o;
  wire n4531_o;
  wire n4532_o;
  wire n4536_o;
  reg [3:0] n4539_o;
  reg [3:0] n4540_o;
  wire [31:0] n4541_o;
  wire [31:0] n4542_o;
  wire [63:0] n4543_o;
  wire n4545_o;
  wire [1:0] n4546_o;
  wire n4552_o;
  wire n4558_o;
  wire n4564_o;
  wire [2:0] n4569_o;
  reg [1:0] n4570_o;
  reg [1:0] n4571_o;
  reg [1:0] n4572_o;
  reg [1:0] n4573_o;
  wire [15:0] n4574_o;
  wire [15:0] n4575_o;
  wire [31:0] n4576_o;
  wire [15:0] n4577_o;
  wire [47:0] n4578_o;
  wire [15:0] n4579_o;
  wire [63:0] n4580_o;
  wire n4582_o;
  wire [2:0] n4583_o;
  wire n4593_o;
  wire n4603_o;
  wire n4613_o;
  wire n4623_o;
  wire n4633_o;
  wire n4643_o;
  wire n4653_o;
  wire [6:0] n4662_o;
  reg n4663_o;
  reg n4664_o;
  reg n4665_o;
  reg n4666_o;
  reg n4667_o;
  reg n4668_o;
  reg n4669_o;
  reg n4670_o;
  wire [7:0] n4671_o;
  wire [7:0] n4672_o;
  wire [15:0] n4673_o;
  wire [7:0] n4674_o;
  wire [23:0] n4675_o;
  wire [7:0] n4676_o;
  wire [31:0] n4677_o;
  wire [7:0] n4678_o;
  wire [39:0] n4679_o;
  wire [7:0] n4680_o;
  wire [47:0] n4681_o;
  wire [7:0] n4682_o;
  wire [55:0] n4683_o;
  wire [7:0] n4684_o;
  wire [63:0] n4685_o;
  wire [7:0] n4686_o;
  wire [7:0] n4688_o;
  wire [63:0] n4689_o;
  wire [7:0] n4690_o;
  wire [7:0] n4691_o;
  wire [63:0] n4692_o;
  wire [7:0] n4693_o;
  wire [7:0] n4694_o;
  wire [63:0] n4695_o;
  wire n4699_o;
  wire n4702_o;
  wire n4703_o;
  wire [31:0] n4704_o;
  wire n4706_o;
  wire [31:0] n4707_o;
  reg [31:0] n4708_o;
  wire n4711_o;
  wire [1:0] n4712_o;
  wire [15:0] n4713_o;
  wire n4715_o;
  wire [15:0] n4716_o;
  wire n4718_o;
  wire [15:0] n4719_o;
  wire n4721_o;
  wire [15:0] n4722_o;
  wire [2:0] n4723_o;
  reg [15:0] n4724_o;
  wire n4727_o;
  wire [2:0] n4728_o;
  wire [7:0] n4729_o;
  wire n4731_o;
  wire [7:0] n4732_o;
  wire n4734_o;
  wire [7:0] n4735_o;
  wire n4737_o;
  wire [7:0] n4738_o;
  wire n4740_o;
  wire [7:0] n4741_o;
  wire n4743_o;
  wire [7:0] n4744_o;
  wire n4746_o;
  wire [7:0] n4747_o;
  wire n4749_o;
  wire [7:0] n4750_o;
  wire [6:0] n4751_o;
  reg [7:0] n4752_o;
  wire [63:0] n4754_o;
  wire [63:0] n4755_o;
  wire [63:0] n4756_o;
  wire [63:0] n4757_o;
  wire [63:0] n4758_o;
  wire [63:0] n4759_o;
  wire [63:0] n4761_o;
  wire n4771_o;
  wire [63:0] altsyncram_i_n4816;
  wire [10:0] n4817_o;
  wire [63:0] altsyncram_i_q_b;
  reg [63:0] n4820_q;
  reg n4821_q;
  reg n4822_q;
  reg n4823_q;
  reg [2:0] n4824_q;
  reg [2:0] n4825_q;
  reg [2:0] n4826_q;
  reg [13:0] n4827_q;
  reg [13:0] n4828_q;
  reg [13:0] n4829_q;
  reg [10:0] n4830_q;
  reg [7:0] n4831_q;
  reg [63:0] n4832_q;
  reg n4833_q;
  reg [63:0] n4834_q;
  reg n4835_q;
  wire [63:0] n4836_o;
  assign dp_readdatavalid_out = dp_readdatavalid_r;
  assign dp_readdata_out = n4836_o;
  /* ../../HW/src/top/sram.vhd:88:8  */
  assign q = altsyncram_i_n4816; // (signal)
  /* ../../HW/src/top/sram.vhd:89:8  */
  assign q_r = n4820_q; // (signal)
  /* ../../HW/src/top/sram.vhd:90:8  */
  assign rden_r = n4821_q; // (signal)
  /* ../../HW/src/top/sram.vhd:91:8  */
  assign rden_rr = n4822_q; // (signal)
  /* ../../HW/src/top/sram.vhd:92:8  */
  assign rden_rrr = n4823_q; // (signal)
  /* ../../HW/src/top/sram.vhd:93:8  */
  assign rd_vector_r = n4824_q; // (signal)
  /* ../../HW/src/top/sram.vhd:94:8  */
  assign rd_vector_rr = n4825_q; // (signal)
  /* ../../HW/src/top/sram.vhd:95:8  */
  assign rd_vector_rrr = n4826_q; // (signal)
  /* ../../HW/src/top/sram.vhd:96:8  */
  assign valid = n4519_o; // (signal)
  /* ../../HW/src/top/sram.vhd:97:8  */
  assign dp_wr_addr = n4526_o; // (signal)
  /* ../../HW/src/top/sram.vhd:99:8  */
  assign rd_addr_r = n4827_q; // (signal)
  /* ../../HW/src/top/sram.vhd:100:8  */
  assign rd_addr_rr = n4828_q; // (signal)
  /* ../../HW/src/top/sram.vhd:101:8  */
  assign rd_addr_rrr = n4829_q; // (signal)
  /* ../../HW/src/top/sram.vhd:102:8  */
  assign byteena = n4694_o; // (signal)
  /* ../../HW/src/top/sram.vhd:103:8  */
  assign dp_writedata = n4695_o; // (signal)
  /* ../../HW/src/top/sram.vhd:104:8  */
  assign wr_addr_r = n4830_q; // (signal)
  /* ../../HW/src/top/sram.vhd:105:8  */
  assign byteena_r = n4831_q; // (signal)
  /* ../../HW/src/top/sram.vhd:106:8  */
  assign writedata_r = n4832_q; // (signal)
  /* ../../HW/src/top/sram.vhd:107:8  */
  assign wren_r = n4833_q; // (signal)
  /* ../../HW/src/top/sram.vhd:108:8  */
  assign dp_readdata_r = n4834_q; // (signal)
  /* ../../HW/src/top/sram.vhd:109:8  */
  assign dp_readdatavalid = delay_i1_n4522; // (signal)
  /* ../../HW/src/top/sram.vhd:110:8  */
  assign dp_readdatavalid_r = n4835_q; // (signal)
  /* ../../HW/src/top/sram.vhd:114:21  */
  assign n4519_o = dp_read_in & dp_read_gen_valid_in;
  /* ../../HW/src/top/sram.vhd:118:86  */
  assign delay_i1_n4522 = delay_i1_out_out; // (signal)
  /* ../../HW/src/top/sram.vhd:117:1  */
  delay_3 delay_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .in_in(valid),
    .enable_in(n4523_o),
    .out_out(delay_i1_out_out));
  /* ../../HW/src/top/sram.vhd:119:28  */
  assign n4526_o = dp_wr_addr_in[13:3];
  /* ../../HW/src/top/sram.vhd:124:32  */
  assign n4531_o = dp_write_vector_in == 3'b011;
  /* ../../HW/src/top/sram.vhd:125:23  */
  assign n4532_o = dp_wr_addr_in[2];
  /* ../../HW/src/top/sram.vhd:126:9  */
  assign n4536_o = n4532_o == 1'b0;
  /* ../../HW/src/top/sram.vhd:125:5  */
  always @*
    case (n4536_o)
      1'b1: n4539_o = 4'b1111;
      default: n4539_o = 4'b0000;
    endcase
  /* ../../HW/src/top/sram.vhd:125:5  */
  always @*
    case (n4536_o)
      1'b1: n4540_o = 4'b0000;
      default: n4540_o = 4'b1111;
    endcase
  /* ../../HW/src/top/sram.vhd:133:36  */
  assign n4541_o = dp_writedata_in[31:0];
  /* ../../HW/src/top/sram.vhd:134:36  */
  assign n4542_o = dp_writedata_in[31:0];
  /* ../../HW/src/top/sram.vhd:133:68  */
  assign n4543_o = {n4541_o, n4542_o};
  /* ../../HW/src/top/sram.vhd:135:35  */
  assign n4545_o = dp_write_vector_in == 3'b001;
  /* ../../HW/src/top/sram.vhd:136:23  */
  assign n4546_o = dp_wr_addr_in[2:1];
  /* ../../HW/src/top/sram.vhd:137:9  */
  assign n4552_o = n4546_o == 2'b00;
  /* ../../HW/src/top/sram.vhd:142:9  */
  assign n4558_o = n4546_o == 2'b01;
  /* ../../HW/src/top/sram.vhd:147:9  */
  assign n4564_o = n4546_o == 2'b10;
  /* ../../HW/src/pcore/core.vhd:330:10  */
  assign n4569_o = {n4564_o, n4558_o, n4552_o};
  /* ../../HW/src/top/sram.vhd:136:5  */
  always @*
    case (n4569_o)
      3'b100: n4570_o = 2'b00;
      3'b010: n4570_o = 2'b00;
      3'b001: n4570_o = 2'b11;
      default: n4570_o = 2'b00;
    endcase
  /* ../../HW/src/top/sram.vhd:136:5  */
  always @*
    case (n4569_o)
      3'b100: n4571_o = 2'b00;
      3'b010: n4571_o = 2'b11;
      3'b001: n4571_o = 2'b00;
      default: n4571_o = 2'b00;
    endcase
  /* ../../HW/src/top/sram.vhd:136:5  */
  always @*
    case (n4569_o)
      3'b100: n4572_o = 2'b11;
      3'b010: n4572_o = 2'b00;
      3'b001: n4572_o = 2'b00;
      default: n4572_o = 2'b00;
    endcase
  /* ../../HW/src/top/sram.vhd:136:5  */
  always @*
    case (n4569_o)
      3'b100: n4573_o = 2'b00;
      3'b010: n4573_o = 2'b00;
      3'b001: n4573_o = 2'b00;
      default: n4573_o = 2'b11;
    endcase
  /* ../../HW/src/top/sram.vhd:158:36  */
  assign n4574_o = dp_writedata_in[15:0];
  /* ../../HW/src/top/sram.vhd:159:36  */
  assign n4575_o = dp_writedata_in[15:0];
  /* ../../HW/src/top/sram.vhd:158:68  */
  assign n4576_o = {n4574_o, n4575_o};
  /* ../../HW/src/top/sram.vhd:160:36  */
  assign n4577_o = dp_writedata_in[15:0];
  /* ../../HW/src/top/sram.vhd:159:68  */
  assign n4578_o = {n4576_o, n4577_o};
  /* ../../HW/src/top/sram.vhd:161:36  */
  assign n4579_o = dp_writedata_in[15:0];
  /* ../../HW/src/top/sram.vhd:160:68  */
  assign n4580_o = {n4578_o, n4579_o};
  /* ../../HW/src/top/sram.vhd:162:35  */
  assign n4582_o = dp_write_vector_in == 3'b000;
  /* ../../HW/src/top/sram.vhd:163:23  */
  assign n4583_o = dp_wr_addr_in[2:0];
  /* ../../HW/src/top/sram.vhd:164:9  */
  assign n4593_o = n4583_o == 3'b000;
  /* ../../HW/src/top/sram.vhd:173:9  */
  assign n4603_o = n4583_o == 3'b001;
  /* ../../HW/src/top/sram.vhd:182:9  */
  assign n4613_o = n4583_o == 3'b010;
  /* ../../HW/src/top/sram.vhd:191:9  */
  assign n4623_o = n4583_o == 3'b011;
  /* ../../HW/src/top/sram.vhd:200:9  */
  assign n4633_o = n4583_o == 3'b100;
  /* ../../HW/src/top/sram.vhd:209:9  */
  assign n4643_o = n4583_o == 3'b101;
  /* ../../HW/src/top/sram.vhd:218:9  */
  assign n4653_o = n4583_o == 3'b110;
  /* ../../HW/src/pcore/core.vhd:312:10  */
  assign n4662_o = {n4653_o, n4643_o, n4633_o, n4623_o, n4613_o, n4603_o, n4593_o};
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4663_o = 1'b0;
      7'b0100000: n4663_o = 1'b0;
      7'b0010000: n4663_o = 1'b0;
      7'b0001000: n4663_o = 1'b0;
      7'b0000100: n4663_o = 1'b0;
      7'b0000010: n4663_o = 1'b0;
      7'b0000001: n4663_o = 1'b1;
      default: n4663_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4664_o = 1'b0;
      7'b0100000: n4664_o = 1'b0;
      7'b0010000: n4664_o = 1'b0;
      7'b0001000: n4664_o = 1'b0;
      7'b0000100: n4664_o = 1'b0;
      7'b0000010: n4664_o = 1'b1;
      7'b0000001: n4664_o = 1'b0;
      default: n4664_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4665_o = 1'b0;
      7'b0100000: n4665_o = 1'b0;
      7'b0010000: n4665_o = 1'b0;
      7'b0001000: n4665_o = 1'b0;
      7'b0000100: n4665_o = 1'b1;
      7'b0000010: n4665_o = 1'b0;
      7'b0000001: n4665_o = 1'b0;
      default: n4665_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4666_o = 1'b0;
      7'b0100000: n4666_o = 1'b0;
      7'b0010000: n4666_o = 1'b0;
      7'b0001000: n4666_o = 1'b1;
      7'b0000100: n4666_o = 1'b0;
      7'b0000010: n4666_o = 1'b0;
      7'b0000001: n4666_o = 1'b0;
      default: n4666_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4667_o = 1'b0;
      7'b0100000: n4667_o = 1'b0;
      7'b0010000: n4667_o = 1'b1;
      7'b0001000: n4667_o = 1'b0;
      7'b0000100: n4667_o = 1'b0;
      7'b0000010: n4667_o = 1'b0;
      7'b0000001: n4667_o = 1'b0;
      default: n4667_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4668_o = 1'b0;
      7'b0100000: n4668_o = 1'b1;
      7'b0010000: n4668_o = 1'b0;
      7'b0001000: n4668_o = 1'b0;
      7'b0000100: n4668_o = 1'b0;
      7'b0000010: n4668_o = 1'b0;
      7'b0000001: n4668_o = 1'b0;
      default: n4668_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4669_o = 1'b1;
      7'b0100000: n4669_o = 1'b0;
      7'b0010000: n4669_o = 1'b0;
      7'b0001000: n4669_o = 1'b0;
      7'b0000100: n4669_o = 1'b0;
      7'b0000010: n4669_o = 1'b0;
      7'b0000001: n4669_o = 1'b0;
      default: n4669_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram.vhd:163:5  */
  always @*
    case (n4662_o)
      7'b1000000: n4670_o = 1'b0;
      7'b0100000: n4670_o = 1'b0;
      7'b0010000: n4670_o = 1'b0;
      7'b0001000: n4670_o = 1'b0;
      7'b0000100: n4670_o = 1'b0;
      7'b0000010: n4670_o = 1'b0;
      7'b0000001: n4670_o = 1'b0;
      default: n4670_o = 1'b1;
    endcase
  /* ../../HW/src/top/sram.vhd:237:36  */
  assign n4671_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:238:36  */
  assign n4672_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:237:68  */
  assign n4673_o = {n4671_o, n4672_o};
  /* ../../HW/src/top/sram.vhd:239:36  */
  assign n4674_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:238:68  */
  assign n4675_o = {n4673_o, n4674_o};
  /* ../../HW/src/top/sram.vhd:240:36  */
  assign n4676_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:239:68  */
  assign n4677_o = {n4675_o, n4676_o};
  /* ../../HW/src/top/sram.vhd:241:36  */
  assign n4678_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:240:68  */
  assign n4679_o = {n4677_o, n4678_o};
  /* ../../HW/src/top/sram.vhd:242:36  */
  assign n4680_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:241:68  */
  assign n4681_o = {n4679_o, n4680_o};
  /* ../../HW/src/top/sram.vhd:243:36  */
  assign n4682_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:242:68  */
  assign n4683_o = {n4681_o, n4682_o};
  /* ../../HW/src/top/sram.vhd:244:36  */
  assign n4684_o = dp_writedata_in[7:0];
  /* ../../HW/src/top/sram.vhd:243:68  */
  assign n4685_o = {n4683_o, n4684_o};
  assign n4686_o = {n4670_o, n4669_o, n4668_o, n4667_o, n4666_o, n4665_o, n4664_o, n4663_o};
  /* ../../HW/src/top/sram.vhd:162:1  */
  assign n4688_o = n4582_o ? n4686_o : 8'b11111111;
  /* ../../HW/src/top/sram.vhd:162:1  */
  assign n4689_o = n4582_o ? n4685_o : dp_writedata_in;
  /* ../../HW/src/pcore/core.vhd:342:10  */
  assign n4690_o = {n4573_o, n4572_o, n4571_o, n4570_o};
  /* ../../HW/src/top/sram.vhd:135:1  */
  assign n4691_o = n4545_o ? n4690_o : n4688_o;
  /* ../../HW/src/top/sram.vhd:135:1  */
  assign n4692_o = n4545_o ? n4580_o : n4689_o;
  assign n4693_o = {n4540_o, n4539_o};
  /* ../../HW/src/top/sram.vhd:124:1  */
  assign n4694_o = n4531_o ? n4693_o : n4691_o;
  /* ../../HW/src/top/sram.vhd:124:1  */
  assign n4695_o = n4531_o ? n4543_o : n4692_o;
  /* ../../HW/src/top/sram.vhd:253:12  */
  assign n4699_o = ~reset_in;
  /* ../../HW/src/top/sram.vhd:260:31  */
  assign n4702_o = rd_vector_rrr == 3'b011;
  /* ../../HW/src/top/sram.vhd:261:25  */
  assign n4703_o = rd_addr_rrr[2];
  /* ../../HW/src/top/sram.vhd:263:68  */
  assign n4704_o = q_r[31:0];
  /* ../../HW/src/top/sram.vhd:262:13  */
  assign n4706_o = n4703_o == 1'b0;
  /* ../../HW/src/top/sram.vhd:265:68  */
  assign n4707_o = q_r[63:32];
  /* ../../HW/src/top/sram.vhd:261:9  */
  always @*
    case (n4706_o)
      1'b1: n4708_o = n4704_o;
      default: n4708_o = n4707_o;
    endcase
  /* ../../HW/src/top/sram.vhd:268:34  */
  assign n4711_o = rd_vector_rrr == 3'b001;
  /* ../../HW/src/top/sram.vhd:269:25  */
  assign n4712_o = rd_addr_rrr[2:1];
  /* ../../HW/src/top/sram.vhd:271:68  */
  assign n4713_o = q_r[15:0];
  /* ../../HW/src/top/sram.vhd:270:13  */
  assign n4715_o = n4712_o == 2'b00;
  /* ../../HW/src/top/sram.vhd:273:68  */
  assign n4716_o = q_r[31:16];
  /* ../../HW/src/top/sram.vhd:272:13  */
  assign n4718_o = n4712_o == 2'b01;
  /* ../../HW/src/top/sram.vhd:275:68  */
  assign n4719_o = q_r[47:32];
  /* ../../HW/src/top/sram.vhd:274:13  */
  assign n4721_o = n4712_o == 2'b10;
  /* ../../HW/src/top/sram.vhd:277:68  */
  assign n4722_o = q_r[63:48];
  /* ../../HW/src/pcore/core.vhd:345:10  */
  assign n4723_o = {n4721_o, n4718_o, n4715_o};
  /* ../../HW/src/top/sram.vhd:269:9  */
  always @*
    case (n4723_o)
      3'b100: n4724_o = n4719_o;
      3'b010: n4724_o = n4716_o;
      3'b001: n4724_o = n4713_o;
      default: n4724_o = n4722_o;
    endcase
  /* ../../HW/src/top/sram.vhd:280:34  */
  assign n4727_o = rd_vector_rrr == 3'b000;
  /* ../../HW/src/top/sram.vhd:281:25  */
  assign n4728_o = rd_addr_rrr[2:0];
  /* ../../HW/src/top/sram.vhd:283:68  */
  assign n4729_o = q_r[7:0];
  /* ../../HW/src/top/sram.vhd:282:13  */
  assign n4731_o = n4728_o == 3'b000;
  /* ../../HW/src/top/sram.vhd:285:68  */
  assign n4732_o = q_r[15:8];
  /* ../../HW/src/top/sram.vhd:284:13  */
  assign n4734_o = n4728_o == 3'b001;
  /* ../../HW/src/top/sram.vhd:287:68  */
  assign n4735_o = q_r[23:16];
  /* ../../HW/src/top/sram.vhd:286:13  */
  assign n4737_o = n4728_o == 3'b010;
  /* ../../HW/src/top/sram.vhd:289:68  */
  assign n4738_o = q_r[31:24];
  /* ../../HW/src/top/sram.vhd:288:13  */
  assign n4740_o = n4728_o == 3'b011;
  /* ../../HW/src/top/sram.vhd:291:68  */
  assign n4741_o = q_r[39:32];
  /* ../../HW/src/top/sram.vhd:290:13  */
  assign n4743_o = n4728_o == 3'b100;
  /* ../../HW/src/top/sram.vhd:293:68  */
  assign n4744_o = q_r[47:40];
  /* ../../HW/src/top/sram.vhd:292:13  */
  assign n4746_o = n4728_o == 3'b101;
  /* ../../HW/src/top/sram.vhd:295:68  */
  assign n4747_o = q_r[55:48];
  /* ../../HW/src/top/sram.vhd:294:13  */
  assign n4749_o = n4728_o == 3'b110;
  /* ../../HW/src/top/sram.vhd:297:68  */
  assign n4750_o = q_r[63:56];
  /* ../../HW/src/pcore/core.vhd:492:5  */
  assign n4751_o = {n4749_o, n4746_o, n4743_o, n4740_o, n4737_o, n4734_o, n4731_o};
  /* ../../HW/src/top/sram.vhd:281:9  */
  always @*
    case (n4751_o)
      7'b1000000: n4752_o = n4747_o;
      7'b0100000: n4752_o = n4744_o;
      7'b0010000: n4752_o = n4741_o;
      7'b0001000: n4752_o = n4738_o;
      7'b0000100: n4752_o = n4735_o;
      7'b0000010: n4752_o = n4732_o;
      7'b0000001: n4752_o = n4729_o;
      default: n4752_o = n4750_o;
    endcase
  /* ../../HW/src/pcore/core.vhd:492:5  */
  assign n4754_o = {56'b00000000000000000000000000000000000000000000000000000000, n4752_o};
  /* ../../HW/src/top/sram.vhd:280:5  */
  assign n4755_o = n4727_o ? n4754_o : q_r;
  /* ../../HW/src/pcore/core.vhd:492:5  */
  assign n4756_o = {48'b000000000000000000000000000000000000000000000000, n4724_o};
  /* ../../HW/src/top/sram.vhd:268:5  */
  assign n4757_o = n4711_o ? n4756_o : n4755_o;
  /* ../../HW/src/pcore/core.vhd:492:5  */
  assign n4758_o = {32'b00000000000000000000000000000000, n4708_o};
  /* ../../HW/src/top/sram.vhd:260:5  */
  assign n4759_o = n4702_o ? n4758_o : n4757_o;
  /* ../../HW/src/top/sram.vhd:259:1  */
  assign n4761_o = rden_rrr ? n4759_o : 64'b0000000000000000000000000000000000000000000000000000000000000000;
  /* ../../HW/src/top/sram.vhd:312:17  */
  assign n4771_o = ~reset_in;
  /* ../../HW/src/top/sram.vhd:364:16  */
  assign altsyncram_i_n4816 = altsyncram_i_q_b; // (signal)
  /* ../../HW/src/top/sram.vhd:363:31  */
  assign n4817_o = rd_addr_r[13:3];
  /* ../../HW/src/top/sram.vhd:348:1  */
  dpram_be_2048_2048_11_11_64_64 altsyncram_i (
    .address_a(wr_addr_r),
    .byteena_a(byteena_r),
    .clock0(clock_in),
    .data_a(writedata_r),
    .wren_a(wren_r),
    .address_b(n4817_o),
    .q_b(altsyncram_i_q_b));
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4820_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n4820_q <= q;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4821_q <= 1'b0;
    else
      n4821_q <= dp_read_in;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4822_q <= 1'b0;
    else
      n4822_q <= rden_r;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4823_q <= 1'b0;
    else
      n4823_q <= rden_rr;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4824_q <= 3'b000;
    else
      n4824_q <= dp_read_vector_in;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4825_q <= 3'b000;
    else
      n4825_q <= rd_vector_r;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4826_q <= 3'b000;
    else
      n4826_q <= rd_vector_rr;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4827_q <= 14'b00000000000000;
    else
      n4827_q <= dp_rd_addr_in;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4828_q <= 14'b00000000000000;
    else
      n4828_q <= rd_addr_r;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4829_q <= 14'b00000000000000;
    else
      n4829_q <= rd_addr_rr;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4830_q <= 11'b00000000000;
    else
      n4830_q <= dp_wr_addr;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4831_q <= 8'b00000000;
    else
      n4831_q <= byteena;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4832_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n4832_q <= dp_writedata;
  /* ../../HW/src/top/sram.vhd:328:9  */
  always @(posedge clock_in or posedge n4771_o)
    if (n4771_o)
      n4833_q <= 1'b0;
    else
      n4833_q <= dp_write_in;
  /* ../../HW/src/top/sram.vhd:257:1  */
  always @(posedge clock_in or posedge n4699_o)
    if (n4699_o)
      n4834_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n4834_q <= n4761_o;
  /* ../../HW/src/top/sram.vhd:257:1  */
  always @(posedge clock_in or posedge n4699_o)
    if (n4699_o)
      n4835_q <= 1'b0;
    else
      n4835_q <= dp_readdatavalid;
  /* ../../HW/src/top/sram.vhd:115:34  */
  assign n4836_o = dp_readdatavalid_r ? dp_readdata_r : 64'bz;
endmodule

module scfifo_32_6_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [31:0] data_in,
   input  write_in,
   input  read_in,
   output [31:0] q_out,
   output [5:0] ravail_out,
   output [5:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [31:0] q;
  wire [5:0] address_a;
  wire [5:0] address_b;
  wire [5:0] waddr_r;
  wire [5:0] waddr_rr;
  wire [5:0] raddr_r;
  wire [5:0] raddr;
  wire [5:0] ravail;
  wire [5:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [31:0] ram_i_n4450;
  wire [31:0] ram_i_q_b;
  wire [5:0] n4453_o;
  wire [5:0] n4454_o;
  wire n4455_o;
  wire n4458_o;
  wire n4459_o;
  wire [5:0] n4462_o;
  wire [5:0] n4463_o;
  wire n4466_o;
  wire [5:0] n4469_o;
  wire [5:0] n4471_o;
  wire n4472_o;
  wire n4475_o;
  wire [5:0] n4477_o;
  wire n4478_o;
  wire n4481_o;
  wire n4483_o;
  wire n4485_o;
  wire n4488_o;
  wire [5:0] n4510_o;
  reg [5:0] n4511_q;
  reg [5:0] n4512_q;
  reg [5:0] n4513_q;
  reg n4515_q;
  reg n4516_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n4455_o;
  assign full_out = full_r;
  assign almost_full_out = n4459_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n4450; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n4511_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n4512_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n4513_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n4463_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n4453_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n4454_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n4515_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n4516_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n4450 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_64_64_6_6_32_32 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n4453_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n4454_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n4455_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n4458_o = $unsigned(wused) >= $unsigned(6'b000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n4459_o = n4458_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n4462_o = raddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n4463_o = read_in ? n4462_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n4466_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n4469_o = waddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n4471_o = waddr_r + 6'b000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n4472_o = n4471_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n4475_o = n4472_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n4477_o = waddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n4478_o = n4477_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n4481_o = n4478_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n4483_o = write_in ? n4475_o : n4481_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n4485_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n4488_o = n4485_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n4510_o = write_in ? n4469_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4466_o)
    if (n4466_o)
      n4511_q <= 6'b000000;
    else
      n4511_q <= n4510_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4466_o)
    if (n4466_o)
      n4512_q <= 6'b000000;
    else
      n4512_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4466_o)
    if (n4466_o)
      n4513_q <= 6'b000000;
    else
      n4513_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4466_o)
    if (n4466_o)
      n4515_q <= 1'b0;
    else
      n4515_q <= n4488_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4466_o)
    if (n4466_o)
      n4516_q <= 1'b0;
    else
      n4516_q <= n4483_o;
endmodule

module scfifo_24_6_1_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clock_in,
   input  reset_in,
   input  [23:0] data_in,
   input  write_in,
   input  read_in,
   output [23:0] q_out,
   output [5:0] ravail_out,
   output [5:0] wused_out,
   output empty_out,
   output full_out,
   output almost_full_out);
  wire [23:0] q;
  wire [5:0] address_a;
  wire [5:0] address_b;
  wire [5:0] waddr_r;
  wire [5:0] waddr_rr;
  wire [5:0] raddr_r;
  wire [5:0] raddr;
  wire [5:0] ravail;
  wire [5:0] wused;
  wire not_empty_r;
  wire full_r;
  wire [23:0] ram_i_n4377;
  wire [23:0] ram_i_q_b;
  wire [5:0] n4380_o;
  wire [5:0] n4381_o;
  wire n4382_o;
  wire n4385_o;
  wire n4386_o;
  wire [5:0] n4389_o;
  wire [5:0] n4390_o;
  wire n4393_o;
  wire [5:0] n4396_o;
  wire [5:0] n4398_o;
  wire n4399_o;
  wire n4402_o;
  wire [5:0] n4404_o;
  wire n4405_o;
  wire n4408_o;
  wire n4410_o;
  wire n4412_o;
  wire n4415_o;
  wire [5:0] n4437_o;
  reg [5:0] n4438_q;
  reg [5:0] n4439_q;
  reg [5:0] n4440_q;
  reg n4442_q;
  reg n4443_q;
  assign q_out = q;
  assign ravail_out = ravail;
  assign wused_out = wused;
  assign empty_out = n4382_o;
  assign full_out = full_r;
  assign almost_full_out = n4386_o;
  /* ../../HW/src/util/fifo.vhd:53:8  */
  assign q = ram_i_n4377; // (signal)
  /* ../../HW/src/util/fifo.vhd:55:8  */
  assign address_a = waddr_r; // (signal)
  /* ../../HW/src/util/fifo.vhd:56:8  */
  assign address_b = raddr; // (signal)
  /* ../../HW/src/util/fifo.vhd:57:8  */
  assign waddr_r = n4438_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:58:8  */
  assign waddr_rr = n4439_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:59:8  */
  assign raddr_r = n4440_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:60:8  */
  assign raddr = n4390_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:62:8  */
  assign ravail = n4380_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:63:8  */
  assign wused = n4381_o; // (signal)
  /* ../../HW/src/util/fifo.vhd:64:8  */
  assign not_empty_r = n4442_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:65:8  */
  assign full_r = n4443_q; // (signal)
  /* ../../HW/src/util/fifo.vhd:88:16  */
  assign ram_i_n4377 = ram_i_q_b; // (signal)
  /* ../../HW/src/util/fifo.vhd:71:1  */
  dpram_64_64_6_6_24_24 ram_i (
    .address_a(address_a),
    .clock(clock_in),
    .data_a(data_in),
    .wren_a(write_in),
    .address_b(address_b),
    .q_b(ram_i_q_b));
  /* ../../HW/src/util/fifo.vhd:91:20  */
  assign n4380_o = waddr_rr - raddr_r;
  /* ../../HW/src/util/fifo.vhd:92:18  */
  assign n4381_o = waddr_r - raddr_r;
  /* ../../HW/src/util/fifo.vhd:93:14  */
  assign n4382_o = ~not_empty_r;
  /* ../../HW/src/util/fifo.vhd:95:36  */
  assign n4385_o = $unsigned(wused) >= $unsigned(6'b000001);
  /* ../../HW/src/util/fifo.vhd:95:24  */
  assign n4386_o = n4385_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:98:18  */
  assign n4389_o = raddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:98:22  */
  assign n4390_o = read_in ? n4389_o : raddr_r;
  /* ../../HW/src/util/fifo.vhd:110:15  */
  assign n4393_o = ~reset_in;
  /* ../../HW/src/util/fifo.vhd:120:32  */
  assign n4396_o = waddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:121:24  */
  assign n4398_o = waddr_r + 6'b000010;
  /* ../../HW/src/util/fifo.vhd:121:27  */
  assign n4399_o = n4398_o == raddr;
  /* ../../HW/src/util/fifo.vhd:121:13  */
  assign n4402_o = n4399_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:127:24  */
  assign n4404_o = waddr_r + 6'b000001;
  /* ../../HW/src/util/fifo.vhd:127:27  */
  assign n4405_o = n4404_o == raddr;
  /* ../../HW/src/util/fifo.vhd:127:13  */
  assign n4408_o = n4405_o ? 1'b1 : 1'b0;
  /* ../../HW/src/util/fifo.vhd:119:10  */
  assign n4410_o = write_in ? n4402_o : n4408_o;
  /* ../../HW/src/util/fifo.vhd:142:20  */
  assign n4412_o = waddr_r == raddr;
  /* ../../HW/src/util/fifo.vhd:142:10  */
  assign n4415_o = n4412_o ? 1'b0 : 1'b1;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  assign n4437_o = write_in ? n4396_o : waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4393_o)
    if (n4393_o)
      n4438_q <= 6'b000000;
    else
      n4438_q <= n4437_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4393_o)
    if (n4393_o)
      n4439_q <= 6'b000000;
    else
      n4439_q <= waddr_r;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4393_o)
    if (n4393_o)
      n4440_q <= 6'b000000;
    else
      n4440_q <= raddr;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4393_o)
    if (n4393_o)
      n4442_q <= 1'b0;
    else
      n4442_q <= n4415_o;
  /* ../../HW/src/util/fifo.vhd:118:7  */
  always @(posedge clock_in or posedge n4393_o)
    if (n4393_o)
      n4443_q <= 1'b0;
    else
      n4443_q <= n4410_o;
endmodule

module core
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [21:0] dp_rd_addr_in,
   input  dp_rd_fork_in,
   input  dp_rd_addr_mode_in,
   input  [21:0] dp_wr_addr_in,
   input  dp_wr_fork_in,
   input  dp_wr_addr_mode_in,
   input  [5:0] dp_wr_mcast_in,
   input  dp_write_in,
   input  [1:0] dp_write_data_flow_in,
   input  [1:0] dp_write_data_type_in,
   input  [1:0] dp_write_data_model_in,
   input  dp_write_gen_valid_in,
   input  [2:0] dp_write_vector_in,
   input  dp_write_stream_in,
   input  [1:0] dp_write_stream_id_in,
   input  [1:0] dp_write_scatter_in,
   input  dp_read_gen_valid_in,
   input  dp_read_in,
   input  [1:0] dp_read_data_flow_in,
   input  dp_read_stream_in,
   input  [1:0] dp_read_stream_id_in,
   input  [1:0] dp_read_data_type_in,
   input  [1:0] dp_read_data_model_in,
   input  [2:0] dp_read_vector_in,
   input  [1:0] dp_read_scatter_in,
   input  [63:0] dp_writedata_in,
   input  [10:0] task_start_addr_in,
   input  task_in,
   input  task_vm_in,
   input  [4:0] task_pcore_in,
   input  task_lockstep_in,
   input  [3:0] task_tid_mask_in,
   input  [27:0] task_iregister_auto_in,
   input  [1:0] task_data_model_in,
   output dp_write_wait_out,
   output dp_read_wait_out,
   output dp_readdatavalid_out,
   output dp_read_gen_valid_out,
   output [63:0] dp_readdata_out,
   output dp_readdata_vm_out,
   output [1:0] busy_out,
   output ready_out);
  wire [2:0] dp_write_vector_r;
  wire [2:0] dp_write_vector_rr;
  wire [2:0] dp_write_vector_rrr;
  wire [2:0] dp_write_vector_rrrr;
  wire [2:0] dp_write_vector_rrrrr;
  wire [1:0] dp_write_scatter_r;
  wire [1:0] dp_write_scatter_rr;
  wire [1:0] dp_write_scatter_rrr;
  wire [1:0] dp_write_scatter_rrrr;
  wire [1:0] dp_write_scatter_rrrrr;
  wire dp_wr_vm_r;
  wire dp_wr_vm_rr;
  wire dp_wr_vm_rrr;
  wire dp_wr_vm_rrrr;
  wire dp_wr_vm_rrrrr;
  wire dp_code_r;
  wire dp_code_rr;
  wire dp_code_rrr;
  wire dp_code_rrrr;
  wire dp_code_rrrrr;
  wire dp_config_r;
  wire dp_config_rr;
  wire dp_config_rrr;
  wire dp_config_rrrr;
  wire dp_config_rrrrr;
  wire [21:0] dp_wr_addr_r;
  wire [21:0] dp_wr_addr_rr;
  wire [21:0] dp_wr_addr_rrr;
  wire [21:0] dp_wr_addr_rrrr;
  wire [21:0] dp_wr_addr_rrrrr;
  wire [21:0] dp_wr_addr_step_r;
  wire [21:0] dp_wr_addr_step_rr;
  wire [21:0] dp_wr_addr_step_rrr;
  wire [21:0] dp_wr_addr_step_rrrr;
  wire [21:0] dp_wr_addr_step_rrrrr;
  wire dp_wr_share_r;
  wire dp_wr_share_rr;
  wire dp_wr_share_rrr;
  wire dp_wr_share_rrrr;
  wire dp_wr_share_rrrrr;
  wire dp_write_r;
  wire dp_write_rr;
  wire dp_write_rrr;
  wire dp_write_rrrr;
  wire dp_write_rrrrr;
  wire dp_write_gen_valid_r;
  wire dp_write_gen_valid_rr;
  wire dp_write_gen_valid_rrr;
  wire dp_write_gen_valid_rrrr;
  wire dp_write_gen_valid_rrrrr;
  reg [5:0] dp_wr_mcast_r;
  reg [5:0] dp_wr_mcast_rr;
  reg [5:0] dp_wr_mcast_rrr;
  reg [5:0] dp_wr_mcast_rrrr;
  reg [5:0] dp_wr_mcast_rrrrr;
  wire [95:0] dp_writedata_r;
  wire [95:0] dp_writedata_rr;
  wire [95:0] dp_writedata_rrr;
  wire [95:0] dp_writedata_rrrr;
  wire [95:0] dp_writedata_rrrrr;
  wire [95:0] writedata2;
  wire [7:0] dp_stream_read_req_r;
  wire [7:0] dp_stream_read_done_r;
  wire [2:0] dp_read_vector_r;
  wire [1:0] dp_read_scatter_r;
  wire [1:0] dp_read_data_flow_r;
  wire [1:0] dp_read_data_flow2_r;
  wire [1:0] dp_read_data_flow2_rr;
  wire [1:0] dp_read_data_flow2_rrr;
  wire [1:0] dp_read_data_flow2_rrrr;
  wire [1:0] dp_read_data_flow2_rrrrr;
  wire [1:0] dp_read_data_type_r;
  wire dp_read_stream_r;
  wire [1:0] dp_read_stream_id_r;
  wire [1:0] dp_read_stream_id2_r;
  wire dp_rd_vm;
  wire dp_wr_vm;
  wire dp_rd_vm_r;
  wire dp_rd_share;
  wire dp_wr_share;
  wire [21:0] dp_rd_addr;
  wire [21:0] dp_rd_addr_step;
  wire [21:0] dp_wr_addr;
  wire [21:0] dp_wr_addr_step;
  wire [21:0] dp_rd_addr2;
  wire [21:0] dp_wr_addr2;
  wire [1:0] busy;
  wire ready;
  wire [1:0] busy_r;
  wire ready_r;
  wire dp_wr_spe;
  wire dp_wr_pcore_program;
  wire [21:0] dp_rd_addr_r;
  wire [21:0] dp_rd_addr_step_r;
  wire dp_rd_share_r;
  wire dp_read_r;
  wire dp_read_gen_valid_r;
  wire [1:0] dp_rd_page2;
  wire [1:0] dp_wr_page2;
  wire [95:0] writedata;
  wire dp_readdatavalid;
  wire [1:0] dp_readdatavalidv;
  wire dp_read_gen_valid;
  wire dp_readdata_vm;
  wire dp_readdata_vm_r;
  wire dp_readdata_vm_rr;
  wire dp_readdata_vm_rrr;
  wire dp_readdata_vm_rrrr;
  wire dp_readdata_vm_rrrrr;
  wire dp_readdata_vm_rrrrrr;
  wire [1:0] dp_read_data_flow;
  wire dp_read_stream;
  wire [1:0] dp_read_stream_id;
  wire [95:0] dp_readdata;
  wire [95:0] dp_readdata2;
  wire dp_readdatavalid2_r;
  wire dp_readdatavalid2_rr;
  wire dp_readdatavalid2_rrr;
  wire dp_readdatavalid2_rrrr;
  wire dp_readdatavalid2_rrrrr;
  wire dp_readdatavalid2_rrrrrr;
  wire dp_read_gen_valid2_r;
  wire dp_read_gen_valid2_rr;
  wire dp_read_gen_valid2_rrr;
  wire dp_read_gen_valid2_rrrr;
  wire dp_read_gen_valid2_rrrrr;
  wire dp_read_gen_valid2_rrrrrr;
  wire dp_read_stream2_r;
  wire dp_read_stream2_rr;
  wire dp_read_stream2_rrr;
  wire dp_read_stream2_rrrr;
  wire dp_read_stream2_rrrrr;
  wire [95:0] dp_readdata2_r;
  wire [95:0] dp_readdata2_rr;
  wire [95:0] dp_readdata2_rrr;
  wire [95:0] dp_readdata2_rrrr;
  wire [95:0] dp_readdata2_rrrrr;
  wire [1:0] stream_read_id;
  wire [95:0] stream_read_input;
  wire [95:0] stream_read_output;
  wire [1:0] stream_write_id;
  wire [95:0] stream_write_input;
  wire [95:0] stream_write_output;
  wire [2:0] dp_read_vector;
  wire [2:0] dp_read_vaddr;
  wire [95:0] \output ;
  wire [63:0] stream_output_r;
  wire spe_wr;
  wire [8:0] spe_addr;
  wire [23:0] spe_data;
  wire dp_core_write;
  wire dp_core_write_wait_r;
  wire dp_core_write_wait;
  wire dp_core_read;
  wire dp_core_read_wait_r;
  wire dp_write_stream_r;
  wire dp_write_stream_rr;
  wire dp_write_stream_rrr;
  wire dp_write_stream_rrrr;
  wire dp_write_stream_rrrrr;
  wire [1:0] dp_write_stream_id_r;
  wire [79:0] instruction_mu;
  wire [31:0] instruction_imu;
  wire instruction_mu_valid;
  wire instruction_imu_valid;
  wire vm;
  wire [1:0] data_model;
  wire [7:0] enable;
  wire [3:0] tid;
  wire tid_valid1;
  wire [3:0] pre_tid;
  wire pre_tid_valid1;
  wire [3:0] pre_pre_tid;
  wire pre_pre_tid_valid1;
  wire pre_pre_vm;
  wire [1:0] pre_pre_data_model;
  wire [27:0] pre_iregister_auto;
  wire [7:0] i_y_neg;
  wire [7:0] i_y_zero;
  wire n3035_o;
  wire [8:0] n3036_o;
  wire [11:0] n3037_o;
  wire [11:0] n3038_o;
  wire [23:0] n3039_o;
  wire [11:0] n3040_o;
  wire [11:0] gen_stream_n1_stream_i_n3041;
  wire [11:0] gen_stream_n1_stream_i_output_out;
  wire [11:0] n3044_o;
  wire [11:0] gen_stream_n2_stream_i_n3045;
  wire [11:0] gen_stream_n2_stream_i_output_out;
  wire [11:0] n3048_o;
  wire [11:0] gen_stream_n3_stream_i_n3049;
  wire [11:0] gen_stream_n3_stream_i_output_out;
  wire [11:0] n3052_o;
  wire [11:0] gen_stream_n4_stream_i_n3053;
  wire [11:0] gen_stream_n4_stream_i_output_out;
  wire [11:0] n3056_o;
  wire [11:0] gen_stream_n5_stream_i_n3057;
  wire [11:0] gen_stream_n5_stream_i_output_out;
  wire [11:0] n3060_o;
  wire [11:0] gen_stream_n6_stream_i_n3061;
  wire [11:0] gen_stream_n6_stream_i_output_out;
  wire [11:0] n3064_o;
  wire [11:0] gen_stream_n7_stream_i_n3065;
  wire [11:0] gen_stream_n7_stream_i_output_out;
  wire [11:0] n3068_o;
  wire [11:0] gen_stream_n8_stream_i_n3069;
  wire [11:0] gen_stream_n8_stream_i_output_out;
  wire [11:0] n3072_o;
  wire [11:0] gen_stream_1_n1_stream_i1_n3073;
  wire [11:0] gen_stream_1_n1_stream_i1_output_out;
  wire [11:0] n3076_o;
  wire [11:0] gen_stream_1_n2_stream_i1_n3077;
  wire [11:0] gen_stream_1_n2_stream_i1_output_out;
  wire [11:0] n3080_o;
  wire [11:0] gen_stream_1_n3_stream_i1_n3081;
  wire [11:0] gen_stream_1_n3_stream_i1_output_out;
  wire [11:0] n3084_o;
  wire [11:0] gen_stream_1_n4_stream_i1_n3085;
  wire [11:0] gen_stream_1_n4_stream_i1_output_out;
  wire [11:0] n3088_o;
  wire [11:0] gen_stream_1_n5_stream_i1_n3089;
  wire [11:0] gen_stream_1_n5_stream_i1_output_out;
  wire [11:0] n3092_o;
  wire [11:0] gen_stream_1_n6_stream_i1_n3093;
  wire [11:0] gen_stream_1_n6_stream_i1_output_out;
  wire [11:0] n3096_o;
  wire [11:0] gen_stream_1_n7_stream_i1_n3097;
  wire [11:0] gen_stream_1_n7_stream_i1_output_out;
  wire [11:0] n3100_o;
  wire [11:0] gen_stream_1_n8_stream_i1_n3101;
  wire [11:0] gen_stream_1_n8_stream_i1_output_out;
  wire n3107_o;
  wire n3109_o;
  wire n3111_o;
  wire n3112_o;
  wire n3114_o;
  wire [95:0] n3115_o;
  wire n3117_o;
  wire n3118_o;
  wire n3119_o;
  wire n3120_o;
  wire n3122_o;
  wire n3123_o;
  wire n3124_o;
  wire n3125_o;
  wire n3126_o;
  wire n3127_o;
  wire n3130_o;
  wire n3133_o;
  wire [11:0] n3135_o;
  wire [7:0] n3141_o;
  wire [11:0] n3144_o;
  wire [7:0] n3150_o;
  wire [11:0] n3153_o;
  wire [7:0] n3159_o;
  wire [11:0] n3162_o;
  wire [7:0] n3168_o;
  wire [11:0] n3171_o;
  wire [7:0] n3177_o;
  wire [11:0] n3180_o;
  wire [7:0] n3186_o;
  wire [11:0] n3189_o;
  wire [7:0] n3195_o;
  wire [11:0] n3198_o;
  wire [7:0] n3204_o;
  wire [11:0] n3206_o;
  wire [15:0] n3207_o;
  wire [11:0] n3208_o;
  wire [15:0] n3209_o;
  wire [11:0] n3210_o;
  wire [15:0] n3211_o;
  wire [11:0] n3212_o;
  wire [15:0] n3213_o;
  wire [63:0] n3214_o;
  wire [63:0] n3215_o;
  wire [63:0] n3216_o;
  wire n3224_o;
  wire n3225_o;
  wire [47:0] n3226_o;
  wire n3228_o;
  wire [47:0] n3229_o;
  reg [47:0] n3230_o;
  wire n3233_o;
  wire [1:0] n3234_o;
  wire [23:0] n3235_o;
  wire n3237_o;
  wire [23:0] n3238_o;
  wire n3240_o;
  wire [23:0] n3241_o;
  wire n3243_o;
  wire [23:0] n3244_o;
  wire [2:0] n3245_o;
  reg [23:0] n3246_o;
  wire [95:0] n3248_o;
  wire [95:0] n3249_o;
  wire [95:0] n3250_o;
  wire [95:0] n3251_o;
  wire n3255_o;
  wire n3257_o;
  wire n3259_o;
  wire [7:0] n3261_o;
  wire n3363_o;
  wire n3365_o;
  wire [7:0] n3367_o;
  wire n3375_o;
  wire n3376_o;
  wire n3377_o;
  wire n3378_o;
  wire [3:0] n3379_o;
  wire [11:0] n3380_o;
  wire [7:0] n3382_o;
  wire n3390_o;
  wire n3391_o;
  wire n3392_o;
  wire n3393_o;
  wire [3:0] n3394_o;
  wire [11:0] n3395_o;
  wire [7:0] n3397_o;
  wire n3405_o;
  wire n3406_o;
  wire n3407_o;
  wire n3408_o;
  wire [3:0] n3409_o;
  wire [11:0] n3410_o;
  wire [7:0] n3412_o;
  wire n3420_o;
  wire n3421_o;
  wire n3422_o;
  wire n3423_o;
  wire [3:0] n3424_o;
  wire [11:0] n3425_o;
  wire [7:0] n3427_o;
  wire n3435_o;
  wire n3436_o;
  wire n3437_o;
  wire n3438_o;
  wire [3:0] n3439_o;
  wire [11:0] n3440_o;
  wire [7:0] n3442_o;
  wire n3450_o;
  wire n3451_o;
  wire n3452_o;
  wire n3453_o;
  wire [3:0] n3454_o;
  wire [11:0] n3455_o;
  wire [7:0] n3457_o;
  wire n3465_o;
  wire n3466_o;
  wire n3467_o;
  wire n3468_o;
  wire [3:0] n3469_o;
  wire [11:0] n3470_o;
  wire [7:0] n3472_o;
  wire n3480_o;
  wire n3481_o;
  wire n3482_o;
  wire n3483_o;
  wire [3:0] n3484_o;
  wire [11:0] n3485_o;
  wire [7:0] n3487_o;
  wire [11:0] n3496_o;
  wire [7:0] n3498_o;
  wire [11:0] n3507_o;
  wire [7:0] n3509_o;
  wire [11:0] n3518_o;
  wire [7:0] n3520_o;
  wire [11:0] n3529_o;
  wire [7:0] n3531_o;
  wire [11:0] n3540_o;
  wire [7:0] n3542_o;
  wire [11:0] n3551_o;
  wire [7:0] n3553_o;
  wire [11:0] n3562_o;
  wire [7:0] n3564_o;
  wire [11:0] n3573_o;
  wire [95:0] n3574_o;
  wire [95:0] n3575_o;
  wire [95:0] n3576_o;
  wire [15:0] n3577_o;
  wire [11:0] n3578_o;
  wire [15:0] n3579_o;
  wire [11:0] n3580_o;
  wire [15:0] n3581_o;
  wire [11:0] n3582_o;
  wire [15:0] n3583_o;
  wire [11:0] n3584_o;
  wire [95:0] n3589_o;
  wire [95:0] n3590_o;
  wire n3595_o;
  wire n3597_o;
  wire [7:0] n3599_o;
  wire n3601_o;
  wire [2:0] n3604_o;
  wire n3606_o;
  wire [10:0] n3607_o;
  wire [31:0] n3609_o;
  wire [31:0] n3610_o;
  wire n3612_o;
  wire [11:0] n3613_o;
  wire [11:0] n3614_o;
  wire [23:0] n3615_o;
  wire [11:0] n3616_o;
  wire [35:0] n3617_o;
  wire [11:0] n3618_o;
  wire [47:0] n3619_o;
  wire [11:0] n3620_o;
  wire [59:0] n3621_o;
  wire [11:0] n3622_o;
  wire [71:0] n3623_o;
  wire [11:0] n3624_o;
  wire [83:0] n3625_o;
  wire [11:0] n3626_o;
  wire [95:0] n3627_o;
  wire n3629_o;
  wire [23:0] n3630_o;
  wire [23:0] n3631_o;
  wire [47:0] n3632_o;
  wire [23:0] n3633_o;
  wire [71:0] n3634_o;
  wire [23:0] n3635_o;
  wire [95:0] n3636_o;
  wire n3638_o;
  wire [47:0] n3639_o;
  wire [47:0] n3640_o;
  wire [95:0] n3641_o;
  wire [95:0] n3642_o;
  wire [95:0] n3643_o;
  wire [95:0] n3644_o;
  wire [2:0] n3646_o;
  wire [1:0] n3648_o;
  wire n3650_o;
  wire n3653_o;
  wire [21:0] n3654_o;
  wire [21:0] n3655_o;
  wire [21:0] n3656_o;
  wire n3658_o;
  wire n3660_o;
  wire n3662_o;
  wire [5:0] n3664_o;
  wire [63:0] n3665_o;
  wire [63:0] n3666_o;
  wire [63:0] n3667_o;
  wire [31:0] n3668_o;
  wire [31:0] n3669_o;
  wire [31:0] n3670_o;
  wire n3672_o;
  wire [1:0] n3674_o;
  wire [2:0] n3676_o;
  wire [1:0] n3678_o;
  wire n3680_o;
  wire n3682_o;
  wire n3685_o;
  wire [2:0] n3686_o;
  wire [2:0] n3687_o;
  wire [18:0] n3688_o;
  wire [18:0] n3689_o;
  wire [18:0] n3690_o;
  wire [21:0] n3691_o;
  wire n3693_o;
  wire n3695_o;
  wire n3697_o;
  wire [5:0] n3699_o;
  wire [95:0] n3700_o;
  wire [95:0] n3701_o;
  wire [95:0] n3702_o;
  wire n3704_o;
  wire [1:0] n3706_o;
  wire [21:0] n3734_o;
  wire [1:0] n3998_o;
  wire [1:0] n3999_o;
  wire n4002_o;
  wire n4003_o;
  wire n4007_o;
  wire n4008_o;
  wire n4012_o;
  wire n4013_o;
  wire n4017_o;
  wire n4018_o;
  wire n4020_o;
  wire n4021_o;
  wire n4025_o;
  wire n4027_o;
  wire [9:0] n4028_o;
  wire [4:0] n4029_o;
  wire [14:0] n4030_o;
  wire [3:0] n4031_o;
  wire [18:0] n4032_o;
  wire [2:0] n4033_o;
  wire [21:0] n4034_o;
  wire [9:0] n4035_o;
  wire [10:0] n4037_o;
  wire [4:0] n4038_o;
  wire [15:0] n4039_o;
  wire [2:0] n4040_o;
  wire [18:0] n4041_o;
  wire [2:0] n4042_o;
  wire [21:0] n4043_o;
  wire [21:0] n4044_o;
  wire [21:0] n4047_o;
  wire [9:0] n4048_o;
  wire [8:0] n4049_o;
  wire [8:0] n4050_o;
  wire [18:0] n4051_o;
  wire [2:0] n4052_o;
  wire [21:0] n4053_o;
  wire [21:0] n4054_o;
  wire [21:0] n4056_o;
  wire n4061_o;
  wire n4063_o;
  wire [9:0] n4064_o;
  wire [4:0] n4065_o;
  wire [14:0] n4066_o;
  wire [3:0] n4067_o;
  wire [18:0] n4068_o;
  wire [2:0] n4069_o;
  wire [21:0] n4070_o;
  wire [9:0] n4071_o;
  wire [10:0] n4073_o;
  wire [4:0] n4074_o;
  wire [15:0] n4075_o;
  wire [2:0] n4076_o;
  wire [18:0] n4077_o;
  wire [2:0] n4078_o;
  wire [21:0] n4079_o;
  wire [21:0] n4080_o;
  wire [21:0] n4083_o;
  wire [9:0] n4084_o;
  wire [8:0] n4085_o;
  wire [8:0] n4086_o;
  wire [18:0] n4087_o;
  wire [2:0] n4088_o;
  wire [21:0] n4089_o;
  wire [21:0] n4090_o;
  wire [21:0] n4092_o;
  wire [1:0] instr_i_n4094;
  wire instr_i_n4095;
  wire [79:0] instr_i_n4096;
  wire [31:0] instr_i_n4097;
  wire instr_i_n4098;
  wire instr_i_n4099;
  wire instr_i_n4100;
  wire [1:0] instr_i_n4101;
  wire [7:0] instr_i_n4102;
  wire [3:0] instr_i_n4103;
  wire instr_i_n4104;
  wire [3:0] instr_i_n4105;
  wire instr_i_n4106;
  wire [3:0] instr_i_n4107;
  wire instr_i_n4108;
  wire instr_i_n4109;
  wire [1:0] instr_i_n4110;
  wire [27:0] instr_i_n4111;
  wire [1:0] instr_i_busy_out;
  wire instr_i_ready_out;
  wire [79:0] instr_i_instruction_mu_out;
  wire [31:0] instr_i_instruction_imu_out;
  wire instr_i_instruction_mu_valid_out;
  wire instr_i_instruction_imu_valid_out;
  wire instr_i_vm_out;
  wire [1:0] instr_i_data_model_out;
  wire [7:0] instr_i_enable_out;
  wire [3:0] instr_i_tid_out;
  wire instr_i_tid_valid1_out;
  wire [3:0] instr_i_pre_tid_out;
  wire instr_i_pre_tid_valid1_out;
  wire [3:0] instr_i_pre_pre_tid_out;
  wire instr_i_pre_pre_tid_valid1_out;
  wire instr_i_pre_pre_vm_out;
  wire [1:0] instr_i_pre_pre_data_model_out;
  wire [27:0] instr_i_pre_iregister_auto_out;
  wire n4148_o;
  wire [95:0] n4149_o;
  localparam n4150_o = 1'b0;
  localparam n4151_o = 1'b0;
  wire [95:0] gen_cell_n1_cell_i_n4152;
  wire gen_cell_n1_cell_i_n4153;
  wire [2:0] gen_cell_n1_cell_i_n4154;
  wire [2:0] gen_cell_n1_cell_i_n4155;
  wire gen_cell_n1_cell_i_n4156;
  wire gen_cell_n1_cell_i_n4157;
  wire [1:0] gen_cell_n1_cell_i_n4158;
  wire gen_cell_n1_cell_i_n4160;
  wire [1:0] gen_cell_n1_cell_i_n4161;
  wire [3:0] n4162_o;
  wire [3:0] gen_cell_n1_cell_i_n4163;
  wire [3:0] gen_cell_n1_cell_i_n4164;
  wire [95:0] gen_cell_n1_cell_i_dp_readdata_out;
  wire gen_cell_n1_cell_i_dp_readdata_vm_out;
  wire [2:0] gen_cell_n1_cell_i_dp_read_vector_out;
  wire [2:0] gen_cell_n1_cell_i_dp_read_vaddr_out;
  wire gen_cell_n1_cell_i_dp_readdata_valid_out;
  wire gen_cell_n1_cell_i_dp_read_gen_valid_out;
  wire [1:0] gen_cell_n1_cell_i_dp_read_data_flow_out;
  wire [1:0] gen_cell_n1_cell_i_dp_read_data_type_out;
  wire gen_cell_n1_cell_i_dp_read_stream_out;
  wire [1:0] gen_cell_n1_cell_i_dp_read_stream_id_out;
  wire [3:0] gen_cell_n1_cell_i_i_y_neg_out;
  wire [3:0] gen_cell_n1_cell_i_i_y_zero_out;
  localparam n4189_o = 1'b0;
  localparam n4190_o = 1'b0;
  wire [95:0] gen_cell_n2_cell_i_n4191;
  wire gen_cell_n2_cell_i_n4192;
  wire [2:0] gen_cell_n2_cell_i_n4193;
  wire [2:0] gen_cell_n2_cell_i_n4194;
  wire gen_cell_n2_cell_i_n4195;
  wire gen_cell_n2_cell_i_n4196;
  wire [1:0] gen_cell_n2_cell_i_n4197;
  wire gen_cell_n2_cell_i_n4199;
  wire [1:0] gen_cell_n2_cell_i_n4200;
  wire [3:0] n4201_o;
  wire [3:0] gen_cell_n2_cell_i_n4202;
  wire [3:0] gen_cell_n2_cell_i_n4203;
  wire [95:0] gen_cell_n2_cell_i_dp_readdata_out;
  wire gen_cell_n2_cell_i_dp_readdata_vm_out;
  wire [2:0] gen_cell_n2_cell_i_dp_read_vector_out;
  wire [2:0] gen_cell_n2_cell_i_dp_read_vaddr_out;
  wire gen_cell_n2_cell_i_dp_readdata_valid_out;
  wire gen_cell_n2_cell_i_dp_read_gen_valid_out;
  wire [1:0] gen_cell_n2_cell_i_dp_read_data_flow_out;
  wire [1:0] gen_cell_n2_cell_i_dp_read_data_type_out;
  wire gen_cell_n2_cell_i_dp_read_stream_out;
  wire [1:0] gen_cell_n2_cell_i_dp_read_stream_id_out;
  wire [3:0] gen_cell_n2_cell_i_i_y_neg_out;
  wire [3:0] gen_cell_n2_cell_i_i_y_zero_out;
  reg [2:0] n4228_q;
  reg [2:0] n4229_q;
  reg [2:0] n4230_q;
  reg [2:0] n4231_q;
  reg [2:0] n4232_q;
  reg [1:0] n4233_q;
  reg [1:0] n4234_q;
  reg [1:0] n4235_q;
  reg [1:0] n4236_q;
  reg [1:0] n4237_q;
  reg n4238_q;
  reg n4239_q;
  reg n4240_q;
  reg n4241_q;
  reg n4242_q;
  reg n4243_q;
  reg n4244_q;
  reg n4245_q;
  reg n4246_q;
  reg n4247_q;
  reg n4248_q;
  reg n4249_q;
  reg n4250_q;
  reg n4251_q;
  reg n4252_q;
  reg [21:0] n4253_q;
  reg [21:0] n4254_q;
  reg [21:0] n4255_q;
  reg [21:0] n4256_q;
  reg [21:0] n4257_q;
  reg [21:0] n4258_q;
  reg [21:0] n4259_q;
  reg [21:0] n4260_q;
  reg [21:0] n4261_q;
  reg [21:0] n4262_q;
  reg n4263_q;
  reg n4264_q;
  reg n4265_q;
  reg n4266_q;
  reg n4267_q;
  reg n4268_q;
  reg n4269_q;
  reg n4270_q;
  reg n4271_q;
  reg n4272_q;
  reg n4273_q;
  reg n4274_q;
  reg n4275_q;
  reg n4276_q;
  reg n4277_q;
  reg [5:0] n4278_q;
  reg [5:0] n4279_q;
  reg [5:0] n4280_q;
  reg [5:0] n4281_q;
  reg [5:0] n4282_q;
  reg [95:0] n4283_q;
  reg [95:0] n4284_q;
  reg [95:0] n4285_q;
  reg [95:0] n4286_q;
  reg [95:0] n4287_q;
  wire [7:0] n4288_o;
  reg [7:0] n4289_q;
  wire [7:0] n4290_o;
  reg [7:0] n4291_q;
  reg [2:0] n4292_q;
  reg [1:0] n4293_q;
  reg [1:0] n4294_q;
  reg [1:0] n4295_q;
  reg [1:0] n4296_q;
  reg [1:0] n4297_q;
  reg [1:0] n4298_q;
  reg [1:0] n4299_q;
  reg [1:0] n4300_q;
  reg n4306_q;
  reg [1:0] n4307_q;
  reg [1:0] n4308_q;
  reg n4309_q;
  reg [1:0] n4310_q;
  reg n4311_q;
  reg [21:0] n4313_q;
  reg [21:0] n4314_q;
  reg n4315_q;
  reg n4316_q;
  reg n4317_q;
  wire [1:0] n4318_o;
  wire n4319_o;
  wire n4320_o;
  reg n4321_q;
  reg n4322_q;
  reg n4323_q;
  reg n4324_q;
  reg n4325_q;
  reg n4326_q;
  wire [1:0] n4327_o;
  wire n4329_o;
  wire [1:0] n4330_o;
  wire [95:0] n4331_o;
  reg n4332_q;
  reg n4333_q;
  reg n4334_q;
  reg n4335_q;
  reg n4336_q;
  reg n4337_q;
  reg n4338_q;
  reg n4339_q;
  reg n4340_q;
  reg n4341_q;
  reg n4342_q;
  reg n4343_q;
  reg n4344_q;
  reg n4345_q;
  reg n4346_q;
  reg n4347_q;
  reg n4348_q;
  reg [95:0] n4350_q;
  reg [95:0] n4351_q;
  reg [95:0] n4352_q;
  reg [95:0] n4353_q;
  reg [95:0] n4354_q;
  wire [95:0] n4356_o;
  wire [95:0] n4357_o;
  wire [2:0] n4358_o;
  wire [2:0] n4359_o;
  reg [63:0] n4360_q;
  reg n4361_q;
  reg n4362_q;
  reg n4363_q;
  reg n4364_q;
  reg n4365_q;
  reg n4366_q;
  reg n4367_q;
  reg [1:0] n4368_q;
  wire [7:0] n4369_o;
  wire [7:0] n4370_o;
  assign dp_write_wait_out = n3114_o;
  assign dp_read_wait_out = dp_core_read_wait_r;
  assign dp_readdatavalid_out = dp_readdatavalid2_rrrrrr;
  assign dp_read_gen_valid_out = dp_read_gen_valid2_rrrrrr;
  assign dp_readdata_out = stream_output_r;
  assign dp_readdata_vm_out = dp_readdata_vm_rrrrrr;
  assign busy_out = busy_r;
  assign ready_out = ready_r;
  /* ../../HW/src/pcore/core.vhd:91:8  */
  assign dp_write_vector_r = n4228_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:92:8  */
  assign dp_write_vector_rr = n4229_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:93:8  */
  assign dp_write_vector_rrr = n4230_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:94:8  */
  assign dp_write_vector_rrrr = n4231_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:95:8  */
  assign dp_write_vector_rrrrr = n4232_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:97:8  */
  assign dp_write_scatter_r = n4233_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:98:8  */
  assign dp_write_scatter_rr = n4234_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:99:8  */
  assign dp_write_scatter_rrr = n4235_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:100:8  */
  assign dp_write_scatter_rrrr = n4236_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:101:8  */
  assign dp_write_scatter_rrrrr = n4237_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:103:8  */
  assign dp_wr_vm_r = n4238_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:104:8  */
  assign dp_wr_vm_rr = n4239_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:105:8  */
  assign dp_wr_vm_rrr = n4240_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:106:8  */
  assign dp_wr_vm_rrrr = n4241_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:107:8  */
  assign dp_wr_vm_rrrrr = n4242_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:109:8  */
  assign dp_code_r = n4243_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:110:8  */
  assign dp_code_rr = n4244_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:111:8  */
  assign dp_code_rrr = n4245_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:112:8  */
  assign dp_code_rrrr = n4246_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:113:8  */
  assign dp_code_rrrrr = n4247_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:115:8  */
  assign dp_config_r = n4248_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:116:8  */
  assign dp_config_rr = n4249_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:117:8  */
  assign dp_config_rrr = n4250_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:118:8  */
  assign dp_config_rrrr = n4251_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:119:8  */
  assign dp_config_rrrrr = n4252_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:121:8  */
  assign dp_wr_addr_r = n4253_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:122:8  */
  assign dp_wr_addr_rr = n4254_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:123:8  */
  assign dp_wr_addr_rrr = n4255_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:124:8  */
  assign dp_wr_addr_rrrr = n4256_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:125:8  */
  assign dp_wr_addr_rrrrr = n4257_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:127:8  */
  assign dp_wr_addr_step_r = n4258_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:128:8  */
  assign dp_wr_addr_step_rr = n4259_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:129:8  */
  assign dp_wr_addr_step_rrr = n4260_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:130:8  */
  assign dp_wr_addr_step_rrrr = n4261_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:131:8  */
  assign dp_wr_addr_step_rrrrr = n4262_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:133:8  */
  assign dp_wr_share_r = n4263_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:134:8  */
  assign dp_wr_share_rr = n4264_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:135:8  */
  assign dp_wr_share_rrr = n4265_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:136:8  */
  assign dp_wr_share_rrrr = n4266_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:137:8  */
  assign dp_wr_share_rrrrr = n4267_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:139:8  */
  assign dp_write_r = n4268_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:140:8  */
  assign dp_write_rr = n4269_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:141:8  */
  assign dp_write_rrr = n4270_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:142:8  */
  assign dp_write_rrrr = n4271_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:143:8  */
  assign dp_write_rrrrr = n4272_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:145:8  */
  assign dp_write_gen_valid_r = n4273_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:146:8  */
  assign dp_write_gen_valid_rr = n4274_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:147:8  */
  assign dp_write_gen_valid_rrr = n4275_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:148:8  */
  assign dp_write_gen_valid_rrrr = n4276_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:149:8  */
  assign dp_write_gen_valid_rrrrr = n4277_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:151:8  */
  always @*
    dp_wr_mcast_r = n4278_q; // (isignal)
  initial
    dp_wr_mcast_r = 6'b111111;
  /* ../../HW/src/pcore/core.vhd:152:8  */
  always @*
    dp_wr_mcast_rr = n4279_q; // (isignal)
  initial
    dp_wr_mcast_rr = 6'b111111;
  /* ../../HW/src/pcore/core.vhd:153:8  */
  always @*
    dp_wr_mcast_rrr = n4280_q; // (isignal)
  initial
    dp_wr_mcast_rrr = 6'b111111;
  /* ../../HW/src/pcore/core.vhd:154:8  */
  always @*
    dp_wr_mcast_rrrr = n4281_q; // (isignal)
  initial
    dp_wr_mcast_rrrr = 6'b111111;
  /* ../../HW/src/pcore/core.vhd:155:8  */
  always @*
    dp_wr_mcast_rrrrr = n4282_q; // (isignal)
  initial
    dp_wr_mcast_rrrrr = 6'b111111;
  /* ../../HW/src/pcore/core.vhd:157:8  */
  assign dp_writedata_r = n4283_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:158:8  */
  assign dp_writedata_rr = n4284_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:159:8  */
  assign dp_writedata_rrr = n4285_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:160:8  */
  assign dp_writedata_rrrr = n4286_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:161:8  */
  assign dp_writedata_rrrrr = n4287_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:163:8  */
  assign writedata2 = n4149_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:165:8  */
  assign dp_stream_read_req_r = n4289_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:166:8  */
  assign dp_stream_read_done_r = n4291_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:168:8  */
  assign dp_read_vector_r = n4292_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:169:8  */
  assign dp_read_scatter_r = n4293_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:170:8  */
  assign dp_read_data_flow_r = n4294_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:171:8  */
  assign dp_read_data_flow2_r = n4295_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:172:8  */
  assign dp_read_data_flow2_rr = n4296_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:173:8  */
  assign dp_read_data_flow2_rrr = n4297_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:174:8  */
  assign dp_read_data_flow2_rrrr = n4298_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:175:8  */
  assign dp_read_data_flow2_rrrrr = n4299_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:176:8  */
  assign dp_read_data_type_r = n4300_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:182:8  */
  assign dp_read_stream_r = n4306_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:183:8  */
  assign dp_read_stream_id_r = n4307_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:184:8  */
  assign dp_read_stream_id2_r = n4308_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:185:8  */
  assign dp_rd_vm = n4020_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:186:8  */
  assign dp_wr_vm = n4021_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:187:8  */
  assign dp_rd_vm_r = n4309_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:188:8  */
  assign dp_rd_share = n4003_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:189:8  */
  assign dp_wr_share = n4018_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:190:8  */
  assign dp_rd_addr = n4090_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:191:8  */
  assign dp_rd_addr_step = n4092_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:192:8  */
  assign dp_wr_addr = n4054_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:193:8  */
  assign dp_wr_addr_step = n4056_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:194:8  */
  assign dp_rd_addr2 = dp_rd_addr_in; // (signal)
  /* ../../HW/src/pcore/core.vhd:195:8  */
  assign dp_wr_addr2 = dp_wr_addr_in; // (signal)
  /* ../../HW/src/pcore/core.vhd:196:8  */
  assign busy = instr_i_n4094; // (signal)
  /* ../../HW/src/pcore/core.vhd:197:8  */
  assign ready = instr_i_n4095; // (signal)
  /* ../../HW/src/pcore/core.vhd:198:8  */
  assign busy_r = n4310_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:199:8  */
  assign ready_r = n4311_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:201:8  */
  assign dp_wr_spe = n4008_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:202:8  */
  assign dp_wr_pcore_program = n4013_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:203:8  */
  assign dp_rd_addr_r = n4313_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:204:8  */
  assign dp_rd_addr_step_r = n4314_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:205:8  */
  assign dp_rd_share_r = n4315_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:206:8  */
  assign dp_read_r = n4316_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:207:8  */
  assign dp_read_gen_valid_r = n4317_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:208:8  */
  assign dp_rd_page2 = n3998_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:209:8  */
  assign dp_wr_page2 = n3999_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:210:8  */
  assign writedata = n3590_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:211:8  */
  assign dp_readdatavalid = n3112_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:212:8  */
  assign dp_readdatavalidv = n4318_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:213:8  */
  assign dp_read_gen_valid = n4319_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:214:8  */
  assign dp_readdata_vm = n4320_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:215:8  */
  assign dp_readdata_vm_r = n4321_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:216:8  */
  assign dp_readdata_vm_rr = n4322_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:217:8  */
  assign dp_readdata_vm_rrr = n4323_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:218:8  */
  assign dp_readdata_vm_rrrr = n4324_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:219:8  */
  assign dp_readdata_vm_rrrrr = n4325_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:220:8  */
  assign dp_readdata_vm_rrrrrr = n4326_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:221:8  */
  assign dp_read_data_flow = n4327_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:223:8  */
  assign dp_read_stream = n4329_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:224:8  */
  assign dp_read_stream_id = n4330_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:225:8  */
  assign dp_readdata = n4331_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:226:8  */
  assign dp_readdata2 = n3251_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:227:8  */
  assign dp_readdatavalid2_r = n4332_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:228:8  */
  assign dp_readdatavalid2_rr = n4333_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:229:8  */
  assign dp_readdatavalid2_rrr = n4334_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:230:8  */
  assign dp_readdatavalid2_rrrr = n4335_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:231:8  */
  assign dp_readdatavalid2_rrrrr = n4336_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:232:8  */
  assign dp_readdatavalid2_rrrrrr = n4337_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:233:8  */
  assign dp_read_gen_valid2_r = n4338_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:234:8  */
  assign dp_read_gen_valid2_rr = n4339_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:235:8  */
  assign dp_read_gen_valid2_rrr = n4340_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:236:8  */
  assign dp_read_gen_valid2_rrrr = n4341_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:237:8  */
  assign dp_read_gen_valid2_rrrrr = n4342_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:238:8  */
  assign dp_read_gen_valid2_rrrrrr = n4343_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:239:8  */
  assign dp_read_stream2_r = n4344_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:240:8  */
  assign dp_read_stream2_rr = n4345_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:241:8  */
  assign dp_read_stream2_rrr = n4346_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:242:8  */
  assign dp_read_stream2_rrrr = n4347_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:243:8  */
  assign dp_read_stream2_rrrrr = n4348_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:245:8  */
  assign dp_readdata2_r = n4350_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:246:8  */
  assign dp_readdata2_rr = n4351_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:247:8  */
  assign dp_readdata2_rrr = n4352_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:248:8  */
  assign dp_readdata2_rrrr = n4353_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:249:8  */
  assign dp_readdata2_rrrrr = n4354_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:252:8  */
  assign stream_read_id = dp_read_stream_id2_r; // (signal)
  /* ../../HW/src/pcore/core.vhd:253:8  */
  assign stream_read_input = dp_readdata2_r; // (signal)
  /* ../../HW/src/pcore/core.vhd:254:8  */
  assign stream_read_output = n4356_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:256:8  */
  assign stream_write_id = dp_write_stream_id_r; // (signal)
  /* ../../HW/src/pcore/core.vhd:257:8  */
  assign stream_write_input = dp_writedata_r; // (signal)
  /* ../../HW/src/pcore/core.vhd:258:8  */
  assign stream_write_output = n4357_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:260:8  */
  assign dp_read_vector = n4358_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:261:8  */
  assign dp_read_vaddr = n4359_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:265:8  */
  assign \output  = n3115_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:266:8  */
  assign stream_output_r = n4360_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:268:8  */
  assign spe_wr = n3035_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:269:8  */
  assign spe_addr = n3036_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:270:8  */
  assign spe_data = n3039_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:272:8  */
  assign dp_core_write = n3125_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:273:8  */
  assign dp_core_write_wait_r = n4361_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:274:8  */
  assign dp_core_write_wait = n3120_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:275:8  */
  assign dp_core_read = n3127_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:276:8  */
  assign dp_core_read_wait_r = n4362_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:278:8  */
  assign dp_write_stream_r = n4363_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:279:8  */
  assign dp_write_stream_rr = n4364_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:280:8  */
  assign dp_write_stream_rrr = n4365_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:281:8  */
  assign dp_write_stream_rrrr = n4366_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:282:8  */
  assign dp_write_stream_rrrrr = n4367_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:283:8  */
  assign dp_write_stream_id_r = n4368_q; // (signal)
  /* ../../HW/src/pcore/core.vhd:288:8  */
  assign instruction_mu = instr_i_n4096; // (signal)
  /* ../../HW/src/pcore/core.vhd:289:8  */
  assign instruction_imu = instr_i_n4097; // (signal)
  /* ../../HW/src/pcore/core.vhd:290:8  */
  assign instruction_mu_valid = instr_i_n4098; // (signal)
  /* ../../HW/src/pcore/core.vhd:291:8  */
  assign instruction_imu_valid = instr_i_n4099; // (signal)
  /* ../../HW/src/pcore/core.vhd:292:8  */
  assign vm = instr_i_n4100; // (signal)
  /* ../../HW/src/pcore/core.vhd:293:8  */
  assign data_model = instr_i_n4101; // (signal)
  /* ../../HW/src/pcore/core.vhd:294:8  */
  assign enable = instr_i_n4102; // (signal)
  /* ../../HW/src/pcore/core.vhd:295:8  */
  assign tid = instr_i_n4103; // (signal)
  /* ../../HW/src/pcore/core.vhd:296:8  */
  assign tid_valid1 = instr_i_n4104; // (signal)
  /* ../../HW/src/pcore/core.vhd:297:8  */
  assign pre_tid = instr_i_n4105; // (signal)
  /* ../../HW/src/pcore/core.vhd:298:8  */
  assign pre_tid_valid1 = instr_i_n4106; // (signal)
  /* ../../HW/src/pcore/core.vhd:299:8  */
  assign pre_pre_tid = instr_i_n4107; // (signal)
  /* ../../HW/src/pcore/core.vhd:300:8  */
  assign pre_pre_tid_valid1 = instr_i_n4108; // (signal)
  /* ../../HW/src/pcore/core.vhd:301:8  */
  assign pre_pre_vm = instr_i_n4109; // (signal)
  /* ../../HW/src/pcore/core.vhd:302:8  */
  assign pre_pre_data_model = instr_i_n4110; // (signal)
  /* ../../HW/src/pcore/core.vhd:303:8  */
  assign pre_iregister_auto = instr_i_n4111; // (signal)
  /* ../../HW/src/pcore/core.vhd:304:8  */
  assign i_y_neg = n4369_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:305:8  */
  assign i_y_zero = n4370_o; // (signal)
  /* ../../HW/src/pcore/core.vhd:353:23  */
  assign n3035_o = dp_write_in & dp_wr_spe;
  /* ../../HW/src/pcore/core.vhd:354:24  */
  assign n3036_o = dp_wr_addr2[9:1];
  /* ../../HW/src/pcore/core.vhd:355:28  */
  assign n3037_o = dp_writedata_in[27:16];
  /* ../../HW/src/pcore/core.vhd:355:103  */
  assign n3038_o = dp_writedata_in[11:0];
  /* ../../HW/src/pcore/core.vhd:355:86  */
  assign n3039_o = {n3037_o, n3038_o};
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3040_o = stream_read_input[11:0];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n1_stream_i_n3041 = gen_stream_n1_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n1_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3040_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n1_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3044_o = stream_read_input[23:12];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n2_stream_i_n3045 = gen_stream_n2_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n2_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3044_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n2_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3048_o = stream_read_input[35:24];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n3_stream_i_n3049 = gen_stream_n3_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n3_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3048_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n3_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3052_o = stream_read_input[47:36];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n4_stream_i_n3053 = gen_stream_n4_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n4_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3052_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n4_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3056_o = stream_read_input[59:48];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n5_stream_i_n3057 = gen_stream_n5_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n5_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3056_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n5_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3060_o = stream_read_input[71:60];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n6_stream_i_n3061 = gen_stream_n6_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n6_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3060_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n6_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3064_o = stream_read_input[83:72];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n7_stream_i_n3065 = gen_stream_n7_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n7_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3064_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n7_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:374:42  */
  assign n3068_o = stream_read_input[95:84];
  /* ../../HW/src/pcore/core.vhd:375:26  */
  assign gen_stream_n8_stream_i_n3069 = gen_stream_n8_stream_i_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:370:1  */
  stream gen_stream_n8_stream_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_read_id),
    .input_in(n3068_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_n8_stream_i_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3072_o = stream_write_input[11:0];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n1_stream_i1_n3073 = gen_stream_1_n1_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n1_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3072_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n1_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3076_o = stream_write_input[23:12];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n2_stream_i1_n3077 = gen_stream_1_n2_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n2_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3076_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n2_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3080_o = stream_write_input[35:24];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n3_stream_i1_n3081 = gen_stream_1_n3_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n3_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3080_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n3_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3084_o = stream_write_input[47:36];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n4_stream_i1_n3085 = gen_stream_1_n4_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n4_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3084_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n4_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3088_o = stream_write_input[59:48];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n5_stream_i1_n3089 = gen_stream_1_n5_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n5_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3088_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n5_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3092_o = stream_write_input[71:60];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n6_stream_i1_n3093 = gen_stream_1_n6_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n6_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3092_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n6_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3096_o = stream_write_input[83:72];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n7_stream_i1_n3097 = gen_stream_1_n7_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n7_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3096_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n7_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:395:43  */
  assign n3100_o = stream_write_input[95:84];
  /* ../../HW/src/pcore/core.vhd:396:26  */
  assign gen_stream_1_n8_stream_i1_n3101 = gen_stream_1_n8_stream_i1_output_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:391:1  */
  stream gen_stream_1_n8_stream_i1 (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .stream_id_in(stream_write_id),
    .input_in(n3100_o),
    .config_in(spe_wr),
    .config_reg_in(spe_addr),
    .config_data_in(spe_data),
    .output_out(gen_stream_1_n8_stream_i1_output_out));
  /* ../../HW/src/pcore/core.vhd:413:46  */
  assign n3107_o = dp_readdatavalidv[0];
  /* ../../HW/src/pcore/core.vhd:413:26  */
  assign n3109_o = 1'b0 | n3107_o;
  /* ../../HW/src/pcore/core.vhd:413:46  */
  assign n3111_o = dp_readdatavalidv[1];
  /* ../../HW/src/pcore/core.vhd:413:26  */
  assign n3112_o = n3109_o | n3111_o;
  /* ../../HW/src/pcore/core.vhd:421:30  */
  assign n3114_o = task_in | dp_core_write_wait;
  /* ../../HW/src/pcore/core.vhd:433:30  */
  assign n3115_o = dp_read_stream2_rrrrr ? stream_read_output : dp_readdata2_rrrrr;
  /* ../../HW/src/pcore/core.vhd:435:84  */
  assign n3117_o = dp_stream_read_req_r != dp_stream_read_done_r;
  /* ../../HW/src/pcore/core.vhd:435:110  */
  assign n3118_o = dp_write_stream_in & n3117_o;
  /* ../../HW/src/pcore/core.vhd:435:58  */
  assign n3119_o = dp_core_write_wait_r | n3118_o;
  /* ../../HW/src/pcore/core.vhd:435:27  */
  assign n3120_o = n3119_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/core.vhd:436:35  */
  assign n3122_o = ~dp_wr_spe;
  /* ../../HW/src/pcore/core.vhd:436:30  */
  assign n3123_o = dp_write_in & n3122_o;
  /* ../../HW/src/pcore/core.vhd:436:55  */
  assign n3124_o = ~dp_core_write_wait;
  /* ../../HW/src/pcore/core.vhd:436:50  */
  assign n3125_o = n3123_o & n3124_o;
  /* ../../HW/src/pcore/core.vhd:437:33  */
  assign n3126_o = ~dp_core_read_wait_r;
  /* ../../HW/src/pcore/core.vhd:437:28  */
  assign n3127_o = dp_read_in & n3126_o;
  /* ../../HW/src/pcore/core.vhd:445:17  */
  assign n3130_o = ~reset_in;
  /* ../../HW/src/pcore/core.vhd:449:40  */
  assign n3133_o = dp_read_data_flow2_rrrrr == 2'b00;
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3135_o = \output [11:0];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3141_o = n3135_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3144_o = \output [23:12];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3150_o = n3144_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3153_o = \output [35:24];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3159_o = n3153_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3162_o = \output [47:36];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3168_o = n3162_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3171_o = \output [59:48];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3177_o = n3171_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3180_o = \output [71:60];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3186_o = n3180_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3189_o = \output [83:72];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3195_o = n3189_o[7:0];
  /* ../../HW/src/pcore/core.vhd:451:98  */
  assign n3198_o = \output [95:84];
  /* ../../HW/src/pcore/core.vhd:347:21  */
  assign n3204_o = n3198_o[7:0];
  /* ../../HW/src/pcore/core.vhd:455:127  */
  assign n3206_o = \output [11:0];
  /* ../../HW/src/pcore/core.vhd:455:107  */
  assign n3207_o = {{4{n3206_o[11]}}, n3206_o}; // sext
  /* ../../HW/src/pcore/core.vhd:455:127  */
  assign n3208_o = \output [23:12];
  /* ../../HW/src/pcore/core.vhd:455:107  */
  assign n3209_o = {{4{n3208_o[11]}}, n3208_o}; // sext
  /* ../../HW/src/pcore/core.vhd:455:127  */
  assign n3210_o = \output [35:24];
  /* ../../HW/src/pcore/core.vhd:455:107  */
  assign n3211_o = {{4{n3210_o[11]}}, n3210_o}; // sext
  /* ../../HW/src/pcore/core.vhd:455:127  */
  assign n3212_o = \output [47:36];
  /* ../../HW/src/pcore/core.vhd:455:107  */
  assign n3213_o = {{4{n3212_o[11]}}, n3212_o}; // sext
  assign n3214_o = {n3213_o, n3211_o, n3209_o, n3207_o};
  assign n3215_o = {n3204_o, n3195_o, n3186_o, n3177_o, n3168_o, n3159_o, n3150_o, n3141_o};
  /* ../../HW/src/pcore/core.vhd:449:13  */
  assign n3216_o = n3133_o ? n3215_o : n3214_o;
  /* ../../HW/src/pcore/core.vhd:464:28  */
  assign n3224_o = dp_read_vector == 3'b011;
  /* ../../HW/src/pcore/core.vhd:465:22  */
  assign n3225_o = dp_read_vaddr[2];
  /* ../../HW/src/pcore/core.vhd:467:68  */
  assign n3226_o = dp_readdata[47:0];
  /* ../../HW/src/pcore/core.vhd:466:7  */
  assign n3228_o = n3225_o == 1'b0;
  /* ../../HW/src/pcore/core.vhd:469:68  */
  assign n3229_o = dp_readdata[95:48];
  /* ../../HW/src/pcore/core.vhd:465:4  */
  always @*
    case (n3228_o)
      1'b1: n3230_o = n3226_o;
      default: n3230_o = n3229_o;
    endcase
  /* ../../HW/src/pcore/core.vhd:472:31  */
  assign n3233_o = dp_read_vector == 3'b001;
  /* ../../HW/src/pcore/core.vhd:473:22  */
  assign n3234_o = dp_read_vaddr[2:1];
  /* ../../HW/src/pcore/core.vhd:475:68  */
  assign n3235_o = dp_readdata[23:0];
  /* ../../HW/src/pcore/core.vhd:474:7  */
  assign n3237_o = n3234_o == 2'b00;
  /* ../../HW/src/pcore/core.vhd:477:68  */
  assign n3238_o = dp_readdata[47:24];
  /* ../../HW/src/pcore/core.vhd:476:7  */
  assign n3240_o = n3234_o == 2'b01;
  /* ../../HW/src/pcore/core.vhd:479:68  */
  assign n3241_o = dp_readdata[71:48];
  /* ../../HW/src/pcore/core.vhd:478:7  */
  assign n3243_o = n3234_o == 2'b10;
  /* ../../HW/src/pcore/core.vhd:481:68  */
  assign n3244_o = dp_readdata[95:72];
  assign n3245_o = {n3243_o, n3240_o, n3237_o};
  /* ../../HW/src/pcore/core.vhd:473:4  */
  always @*
    case (n3245_o)
      3'b100: n3246_o = n3241_o;
      3'b010: n3246_o = n3238_o;
      3'b001: n3246_o = n3235_o;
      default: n3246_o = n3244_o;
    endcase
  assign n3248_o = {72'b000000000000000000000000000000000000000000000000000000000000000000000000, n3246_o};
  /* ../../HW/src/pcore/core.vhd:472:1  */
  assign n3249_o = n3233_o ? n3248_o : dp_readdata;
  assign n3250_o = {48'b000000000000000000000000000000000000000000000000, n3230_o};
  /* ../../HW/src/pcore/core.vhd:464:1  */
  assign n3251_o = n3224_o ? n3250_o : n3249_o;
  /* ../../HW/src/pcore/core.vhd:492:17  */
  assign n3255_o = ~reset_in;
  /* ../../HW/src/pcore/core.vhd:532:35  */
  assign n3257_o = dp_read_gen_valid & dp_readdatavalid;
  /* ../../HW/src/pcore/core.vhd:532:11  */
  assign n3259_o = n3257_o ? dp_read_stream : 1'b0;
  /* ../../HW/src/pcore/core.vhd:540:60  */
  assign n3261_o = dp_stream_read_done_r + 8'b00000001;
  /* ../../HW/src/pcore/core.vhd:587:25  */
  assign n3363_o = dp_write_data_flow_in == 2'b00;
  /* ../../HW/src/pcore/core.vhd:589:28  */
  assign n3365_o = dp_write_data_type_in == 2'b01;
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3367_o = dp_writedata_in[7:0];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3375_o = n3367_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3376_o = n3367_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3377_o = n3367_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3378_o = n3367_o[7];
  assign n3379_o = {n3375_o, n3376_o, n3377_o, n3378_o};
  assign n3380_o = {n3379_o, n3367_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3382_o = dp_writedata_in[15:8];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3390_o = n3382_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3391_o = n3382_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3392_o = n3382_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3393_o = n3382_o[7];
  assign n3394_o = {n3390_o, n3391_o, n3392_o, n3393_o};
  assign n3395_o = {n3394_o, n3382_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3397_o = dp_writedata_in[23:16];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3405_o = n3397_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3406_o = n3397_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3407_o = n3397_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3408_o = n3397_o[7];
  assign n3409_o = {n3405_o, n3406_o, n3407_o, n3408_o};
  assign n3410_o = {n3409_o, n3397_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3412_o = dp_writedata_in[31:24];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3420_o = n3412_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3421_o = n3412_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3422_o = n3412_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3423_o = n3412_o[7];
  assign n3424_o = {n3420_o, n3421_o, n3422_o, n3423_o};
  assign n3425_o = {n3424_o, n3412_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3427_o = dp_writedata_in[39:32];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3435_o = n3427_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3436_o = n3427_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3437_o = n3427_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3438_o = n3427_o[7];
  assign n3439_o = {n3435_o, n3436_o, n3437_o, n3438_o};
  assign n3440_o = {n3439_o, n3427_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3442_o = dp_writedata_in[47:40];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3450_o = n3442_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3451_o = n3442_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3452_o = n3442_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3453_o = n3442_o[7];
  assign n3454_o = {n3450_o, n3451_o, n3452_o, n3453_o};
  assign n3455_o = {n3454_o, n3442_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3457_o = dp_writedata_in[55:48];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3465_o = n3457_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3466_o = n3457_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3467_o = n3457_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3468_o = n3457_o[7];
  assign n3469_o = {n3465_o, n3466_o, n3467_o, n3468_o};
  assign n3470_o = {n3469_o, n3457_o};
  /* ../../HW/src/pcore/core.vhd:591:100  */
  assign n3472_o = dp_writedata_in[63:56];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3480_o = n3472_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3481_o = n3472_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3482_o = n3472_o[7];
  /* ../../HW/src/pcore/core.vhd:318:70  */
  assign n3483_o = n3472_o[7];
  assign n3484_o = {n3480_o, n3481_o, n3482_o, n3483_o};
  assign n3485_o = {n3484_o, n3472_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3487_o = dp_writedata_in[7:0];
  assign n3496_o = {4'b0000, n3487_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3498_o = dp_writedata_in[15:8];
  assign n3507_o = {4'b0000, n3498_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3509_o = dp_writedata_in[23:16];
  assign n3518_o = {4'b0000, n3509_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3520_o = dp_writedata_in[31:24];
  assign n3529_o = {4'b0000, n3520_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3531_o = dp_writedata_in[39:32];
  assign n3540_o = {4'b0000, n3531_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3542_o = dp_writedata_in[47:40];
  assign n3551_o = {4'b0000, n3542_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3553_o = dp_writedata_in[55:48];
  assign n3562_o = {4'b0000, n3553_o};
  /* ../../HW/src/pcore/core.vhd:595:101  */
  assign n3564_o = dp_writedata_in[63:56];
  assign n3573_o = {4'b0000, n3564_o};
  assign n3574_o = {n3573_o, n3562_o, n3551_o, n3540_o, n3529_o, n3518_o, n3507_o, n3496_o};
  assign n3575_o = {n3485_o, n3470_o, n3455_o, n3440_o, n3425_o, n3410_o, n3395_o, n3380_o};
  /* ../../HW/src/pcore/core.vhd:589:4  */
  assign n3576_o = n3365_o ? n3575_o : n3574_o;
  /* ../../HW/src/pcore/core.vhd:601:117  */
  assign n3577_o = dp_writedata_in[15:0];
  /* ../../HW/src/pcore/core.vhd:601:88  */
  assign n3578_o = n3577_o[11:0];  // trunc
  /* ../../HW/src/pcore/core.vhd:601:117  */
  assign n3579_o = dp_writedata_in[31:16];
  /* ../../HW/src/pcore/core.vhd:601:88  */
  assign n3580_o = n3579_o[11:0];  // trunc
  /* ../../HW/src/pcore/core.vhd:601:117  */
  assign n3581_o = dp_writedata_in[47:32];
  /* ../../HW/src/pcore/core.vhd:601:88  */
  assign n3582_o = n3581_o[11:0];  // trunc
  /* ../../HW/src/pcore/core.vhd:601:117  */
  assign n3583_o = dp_writedata_in[63:48];
  /* ../../HW/src/pcore/core.vhd:601:88  */
  assign n3584_o = n3583_o[11:0];  // trunc
  assign n3589_o = {12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, n3584_o, n3582_o, n3580_o, n3578_o};
  /* ../../HW/src/pcore/core.vhd:587:1  */
  assign n3590_o = n3363_o ? n3576_o : n3589_o;
  /* ../../HW/src/pcore/core.vhd:617:17  */
  assign n3595_o = ~reset_in;
  /* ../../HW/src/pcore/core.vhd:741:33  */
  assign n3597_o = dp_read_stream_in & dp_core_read;
  /* ../../HW/src/pcore/core.vhd:742:61  */
  assign n3599_o = dp_stream_read_req_r + 8'b00000001;
  /* ../../HW/src/pcore/core.vhd:772:30  */
  assign n3601_o = ~task_vm_in;
  /* ../../HW/src/pcore/core.vhd:772:17  */
  assign n3604_o = n3601_o ? 3'b000 : 3'b001;
  /* ../../HW/src/pcore/core.vhd:800:35  */
  assign n3606_o = dp_wr_pcore_program & dp_write_in;
  /* ../../HW/src/pcore/core.vhd:804:78  */
  assign n3607_o = dp_wr_addr_in[12:2];
  /* ../../HW/src/pcore/core.vhd:806:75  */
  assign n3609_o = dp_writedata_in[63:32];
  /* ../../HW/src/pcore/core.vhd:807:88  */
  assign n3610_o = dp_writedata_in[31:0];
  /* ../../HW/src/pcore/core.vhd:828:48  */
  assign n3612_o = dp_write_vector_in == 3'b000;
  /* ../../HW/src/pcore/core.vhd:829:47  */
  assign n3613_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:830:47  */
  assign n3614_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:829:77  */
  assign n3615_o = {n3613_o, n3614_o};
  /* ../../HW/src/pcore/core.vhd:831:47  */
  assign n3616_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:830:77  */
  assign n3617_o = {n3615_o, n3616_o};
  /* ../../HW/src/pcore/core.vhd:832:47  */
  assign n3618_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:831:77  */
  assign n3619_o = {n3617_o, n3618_o};
  /* ../../HW/src/pcore/core.vhd:833:47  */
  assign n3620_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:832:77  */
  assign n3621_o = {n3619_o, n3620_o};
  /* ../../HW/src/pcore/core.vhd:834:47  */
  assign n3622_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:833:77  */
  assign n3623_o = {n3621_o, n3622_o};
  /* ../../HW/src/pcore/core.vhd:835:47  */
  assign n3624_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:834:77  */
  assign n3625_o = {n3623_o, n3624_o};
  /* ../../HW/src/pcore/core.vhd:836:47  */
  assign n3626_o = writedata[11:0];
  /* ../../HW/src/pcore/core.vhd:835:77  */
  assign n3627_o = {n3625_o, n3626_o};
  /* ../../HW/src/pcore/core.vhd:837:51  */
  assign n3629_o = dp_write_vector_in == 3'b001;
  /* ../../HW/src/pcore/core.vhd:838:47  */
  assign n3630_o = writedata[23:0];
  /* ../../HW/src/pcore/core.vhd:839:47  */
  assign n3631_o = writedata[23:0];
  /* ../../HW/src/pcore/core.vhd:838:79  */
  assign n3632_o = {n3630_o, n3631_o};
  /* ../../HW/src/pcore/core.vhd:840:47  */
  assign n3633_o = writedata[23:0];
  /* ../../HW/src/pcore/core.vhd:839:79  */
  assign n3634_o = {n3632_o, n3633_o};
  /* ../../HW/src/pcore/core.vhd:841:47  */
  assign n3635_o = writedata[23:0];
  /* ../../HW/src/pcore/core.vhd:840:79  */
  assign n3636_o = {n3634_o, n3635_o};
  /* ../../HW/src/pcore/core.vhd:842:51  */
  assign n3638_o = dp_write_vector_in == 3'b011;
  /* ../../HW/src/pcore/core.vhd:843:47  */
  assign n3639_o = writedata[47:0];
  /* ../../HW/src/pcore/core.vhd:844:47  */
  assign n3640_o = writedata[47:0];
  /* ../../HW/src/pcore/core.vhd:843:79  */
  assign n3641_o = {n3639_o, n3640_o};
  /* ../../HW/src/pcore/core.vhd:842:17  */
  assign n3642_o = n3638_o ? n3641_o : writedata;
  /* ../../HW/src/pcore/core.vhd:837:17  */
  assign n3643_o = n3629_o ? n3636_o : n3642_o;
  /* ../../HW/src/pcore/core.vhd:828:17  */
  assign n3644_o = n3612_o ? n3627_o : n3643_o;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3646_o = n3606_o ? 3'b000 : dp_write_vector_in;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3648_o = n3606_o ? 2'b00 : dp_write_scatter_in;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3650_o = n3606_o ? 1'b0 : dp_wr_vm;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3653_o = n3606_o ? 1'b1 : 1'b0;
  assign n3654_o = {11'b00000000000, n3607_o};
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3655_o = n3606_o ? n3654_o : dp_wr_addr;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3656_o = n3606_o ? dp_wr_addr_step_r : dp_wr_addr_step;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3658_o = n3606_o ? 1'b0 : dp_wr_share;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3660_o = n3606_o ? 1'b1 : dp_core_write;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3662_o = n3606_o ? 1'b0 : dp_write_gen_valid_in;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3664_o = n3606_o ? 6'b111111 : dp_wr_mcast_in;
  assign n3665_o = {n3610_o, n3609_o};
  assign n3666_o = n3644_o[63:0];
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3667_o = n3606_o ? n3665_o : n3666_o;
  assign n3668_o = n3644_o[95:64];
  assign n3669_o = dp_writedata_r[95:64];
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3670_o = n3606_o ? n3669_o : n3668_o;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3672_o = n3606_o ? 1'b0 : dp_write_stream_in;
  /* ../../HW/src/pcore/core.vhd:800:13  */
  assign n3674_o = n3606_o ? 2'b00 : dp_write_stream_id_in;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3676_o = task_in ? 3'b000 : n3646_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3678_o = task_in ? 2'b00 : n3648_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3680_o = task_in ? 1'b0 : n3650_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3682_o = task_in ? 1'b0 : n3653_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3685_o = task_in ? 1'b1 : 1'b0;
  assign n3686_o = n3655_o[2:0];
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3687_o = task_in ? n3604_o : n3686_o;
  assign n3688_o = n3655_o[21:3];
  assign n3689_o = dp_wr_addr_r[21:3];
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3690_o = task_in ? n3689_o : n3688_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3691_o = task_in ? dp_wr_addr_step_r : n3656_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3693_o = task_in ? 1'b0 : n3658_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3695_o = task_in ? 1'b1 : n3660_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3697_o = task_in ? 1'b0 : n3662_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3699_o = task_in ? 6'b111111 : n3664_o;
  assign n3700_o = {n3670_o, n3667_o};
  assign n3701_o = {45'b000000000000000000000000000000000000000000000, task_data_model_in, task_iregister_auto_in, task_tid_mask_in, task_lockstep_in, task_pcore_in, task_start_addr_in};
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3702_o = task_in ? n3701_o : n3700_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3704_o = task_in ? 1'b0 : n3672_o;
  /* ../../HW/src/pcore/core.vhd:767:13  */
  assign n3706_o = task_in ? 2'b00 : n3674_o;
  assign n3734_o = {n3690_o, n3687_o};
  /* ../../HW/src/pcore/core.vhd:930:36  */
  assign n3998_o = dp_rd_addr2[20:19];
  /* ../../HW/src/pcore/core.vhd:932:36  */
  assign n3999_o = dp_wr_addr2[20:19];
  /* ../../HW/src/pcore/core.vhd:934:37  */
  assign n4002_o = dp_rd_page2 == 2'b00;
  /* ../../HW/src/pcore/core.vhd:934:20  */
  assign n4003_o = n4002_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/core.vhd:936:35  */
  assign n4007_o = dp_wr_page2 == 2'b10;
  /* ../../HW/src/pcore/core.vhd:936:18  */
  assign n4008_o = n4007_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/core.vhd:938:45  */
  assign n4012_o = dp_wr_page2 == 2'b11;
  /* ../../HW/src/pcore/core.vhd:938:28  */
  assign n4013_o = n4012_o ? 1'b1 : 1'b0;
  /* ../../HW/src/pcore/core.vhd:940:37  */
  assign n4017_o = dp_wr_page2 == 2'b00;
  /* ../../HW/src/pcore/core.vhd:940:20  */
  assign n4018_o = n4017_o ? 1'b0 : 1'b1;
  /* ../../HW/src/pcore/core.vhd:942:24  */
  assign n4020_o = dp_rd_addr2[21];
  /* ../../HW/src/pcore/core.vhd:944:24  */
  assign n4021_o = dp_wr_addr2[21];
  /* ../../HW/src/pcore/core.vhd:952:16  */
  assign n4025_o = dp_wr_page2 == 2'b00;
  /* ../../HW/src/pcore/core.vhd:953:29  */
  assign n4027_o = dp_write_data_model_in == 2'b00;
  /* ../../HW/src/pcore/core.vhd:954:32  */
  assign n4028_o = dp_wr_addr2[21:12];
  /* ../../HW/src/pcore/core.vhd:955:32  */
  assign n4029_o = dp_wr_addr2[7:3];
  /* ../../HW/src/pcore/core.vhd:954:91  */
  assign n4030_o = {n4028_o, n4029_o};
  /* ../../HW/src/pcore/core.vhd:956:32  */
  assign n4031_o = dp_wr_addr2[11:8];
  /* ../../HW/src/pcore/core.vhd:955:75  */
  assign n4032_o = {n4030_o, n4031_o};
  /* ../../HW/src/pcore/core.vhd:957:32  */
  assign n4033_o = dp_wr_addr2[2:0];
  /* ../../HW/src/pcore/core.vhd:956:90  */
  assign n4034_o = {n4032_o, n4033_o};
  /* ../../HW/src/pcore/core.vhd:960:32  */
  assign n4035_o = dp_wr_addr2[21:12];
  /* ../../HW/src/pcore/core.vhd:960:91  */
  assign n4037_o = {n4035_o, 1'b0};
  /* ../../HW/src/pcore/core.vhd:962:32  */
  assign n4038_o = dp_wr_addr2[7:3];
  /* ../../HW/src/pcore/core.vhd:961:25  */
  assign n4039_o = {n4037_o, n4038_o};
  /* ../../HW/src/pcore/core.vhd:963:32  */
  assign n4040_o = dp_wr_addr2[10:8];
  /* ../../HW/src/pcore/core.vhd:962:75  */
  assign n4041_o = {n4039_o, n4040_o};
  /* ../../HW/src/pcore/core.vhd:964:32  */
  assign n4042_o = dp_wr_addr2[2:0];
  /* ../../HW/src/pcore/core.vhd:963:92  */
  assign n4043_o = {n4041_o, n4042_o};
  /* ../../HW/src/pcore/core.vhd:953:4  */
  assign n4044_o = n4027_o ? n4034_o : n4043_o;
  /* ../../HW/src/pcore/core.vhd:953:4  */
  assign n4047_o = n4027_o ? 22'b0000000000000010000000 : 22'b0000000000000001000000;
  /* ../../HW/src/pcore/core.vhd:968:29  */
  assign n4048_o = dp_wr_addr2[21:12];
  /* ../../HW/src/pcore/core.vhd:969:33  */
  assign n4049_o = dp_wr_addr2[11:3];
  /* ../../HW/src/pcore/core.vhd:969:18  */
  assign n4050_o = ~n4049_o;
  /* ../../HW/src/pcore/core.vhd:968:88  */
  assign n4051_o = {n4048_o, n4050_o};
  /* ../../HW/src/pcore/core.vhd:970:29  */
  assign n4052_o = dp_wr_addr2[2:0];
  /* ../../HW/src/pcore/core.vhd:969:90  */
  assign n4053_o = {n4051_o, n4052_o};
  /* ../../HW/src/pcore/core.vhd:952:1  */
  assign n4054_o = n4025_o ? n4044_o : n4053_o;
  /* ../../HW/src/pcore/core.vhd:952:1  */
  assign n4056_o = n4025_o ? n4047_o : 22'b0000000000000000000000;
  /* ../../HW/src/pcore/core.vhd:981:16  */
  assign n4061_o = dp_rd_page2 == 2'b00;
  /* ../../HW/src/pcore/core.vhd:982:28  */
  assign n4063_o = dp_read_data_model_in == 2'b00;
  /* ../../HW/src/pcore/core.vhd:983:32  */
  assign n4064_o = dp_rd_addr2[21:12];
  /* ../../HW/src/pcore/core.vhd:984:32  */
  assign n4065_o = dp_rd_addr2[7:3];
  /* ../../HW/src/pcore/core.vhd:983:91  */
  assign n4066_o = {n4064_o, n4065_o};
  /* ../../HW/src/pcore/core.vhd:985:32  */
  assign n4067_o = dp_rd_addr2[11:8];
  /* ../../HW/src/pcore/core.vhd:984:75  */
  assign n4068_o = {n4066_o, n4067_o};
  /* ../../HW/src/pcore/core.vhd:986:32  */
  assign n4069_o = dp_rd_addr2[2:0];
  /* ../../HW/src/pcore/core.vhd:985:90  */
  assign n4070_o = {n4068_o, n4069_o};
  /* ../../HW/src/pcore/core.vhd:989:32  */
  assign n4071_o = dp_rd_addr2[21:12];
  /* ../../HW/src/pcore/core.vhd:989:91  */
  assign n4073_o = {n4071_o, 1'b0};
  /* ../../HW/src/pcore/core.vhd:991:32  */
  assign n4074_o = dp_rd_addr2[7:3];
  /* ../../HW/src/pcore/core.vhd:990:25  */
  assign n4075_o = {n4073_o, n4074_o};
  /* ../../HW/src/pcore/core.vhd:992:32  */
  assign n4076_o = dp_rd_addr2[10:8];
  /* ../../HW/src/pcore/core.vhd:991:75  */
  assign n4077_o = {n4075_o, n4076_o};
  /* ../../HW/src/pcore/core.vhd:993:32  */
  assign n4078_o = dp_rd_addr2[2:0];
  /* ../../HW/src/pcore/core.vhd:992:92  */
  assign n4079_o = {n4077_o, n4078_o};
  /* ../../HW/src/pcore/core.vhd:982:4  */
  assign n4080_o = n4063_o ? n4070_o : n4079_o;
  /* ../../HW/src/pcore/core.vhd:982:4  */
  assign n4083_o = n4063_o ? 22'b0000000000000010000000 : 22'b0000000000000001000000;
  /* ../../HW/src/pcore/core.vhd:997:29  */
  assign n4084_o = dp_rd_addr2[21:12];
  /* ../../HW/src/pcore/core.vhd:998:34  */
  assign n4085_o = dp_rd_addr2[11:3];
  /* ../../HW/src/pcore/core.vhd:998:19  */
  assign n4086_o = ~n4085_o;
  /* ../../HW/src/pcore/core.vhd:997:88  */
  assign n4087_o = {n4084_o, n4086_o};
  /* ../../HW/src/pcore/core.vhd:999:15  */
  assign n4088_o = dp_rd_addr2[2:0];
  /* ../../HW/src/pcore/core.vhd:998:91  */
  assign n4089_o = {n4087_o, n4088_o};
  /* ../../HW/src/pcore/core.vhd:981:1  */
  assign n4090_o = n4061_o ? n4080_o : n4089_o;
  /* ../../HW/src/pcore/core.vhd:981:1  */
  assign n4092_o = n4061_o ? n4083_o : 22'b0000000000000000000000;
  /* ../../HW/src/pcore/core.vhd:1023:25  */
  assign instr_i_n4094 = instr_i_busy_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1024:26  */
  assign instr_i_n4095 = instr_i_ready_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1027:35  */
  assign instr_i_n4096 = instr_i_instruction_mu_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1028:36  */
  assign instr_i_n4097 = instr_i_instruction_imu_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1029:41  */
  assign instr_i_n4098 = instr_i_instruction_mu_valid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1030:42  */
  assign instr_i_n4099 = instr_i_instruction_imu_valid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1031:23  */
  assign instr_i_n4100 = instr_i_vm_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1032:31  */
  assign instr_i_n4101 = instr_i_data_model_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1033:27  */
  assign instr_i_n4102 = instr_i_enable_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1034:24  */
  assign instr_i_n4103 = instr_i_tid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1035:31  */
  assign instr_i_n4104 = instr_i_tid_valid1_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1036:29  */
  assign instr_i_n4105 = instr_i_pre_tid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1037:35  */
  assign instr_i_n4106 = instr_i_pre_tid_valid1_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1038:32  */
  assign instr_i_n4107 = instr_i_pre_pre_tid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1039:39  */
  assign instr_i_n4108 = instr_i_pre_pre_tid_valid1_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1040:31  */
  assign instr_i_n4109 = instr_i_pre_pre_vm_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1041:39  */
  assign instr_i_n4110 = instr_i_pre_pre_data_model_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1042:39  */
  assign instr_i_n4111 = instr_i_pre_iregister_auto_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1008:1  */
  instr instr_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .dp_code_in(dp_code_r),
    .dp_config_in(dp_config_r),
    .dp_wr_addr_in(dp_wr_addr_r),
    .dp_write_in(dp_write_r),
    .dp_writedata_in(dp_writedata_r),
    .i_y_neg_in(i_y_neg),
    .i_y_zero_in(i_y_zero),
    .busy_out(instr_i_busy_out),
    .ready_out(instr_i_ready_out),
    .instruction_mu_out(instr_i_instruction_mu_out),
    .instruction_imu_out(instr_i_instruction_imu_out),
    .instruction_mu_valid_out(instr_i_instruction_mu_valid_out),
    .instruction_imu_valid_out(instr_i_instruction_imu_valid_out),
    .vm_out(instr_i_vm_out),
    .data_model_out(instr_i_data_model_out),
    .enable_out(instr_i_enable_out),
    .tid_out(instr_i_tid_out),
    .tid_valid1_out(instr_i_tid_valid1_out),
    .pre_tid_out(instr_i_pre_tid_out),
    .pre_tid_valid1_out(instr_i_pre_tid_valid1_out),
    .pre_pre_tid_out(instr_i_pre_pre_tid_out),
    .pre_pre_tid_valid1_out(instr_i_pre_pre_tid_valid1_out),
    .pre_pre_vm_out(instr_i_pre_pre_vm_out),
    .pre_pre_data_model_out(instr_i_pre_pre_data_model_out),
    .pre_iregister_auto_out(instr_i_pre_iregister_auto_out));
  /* ../../HW/src/pcore/core.vhd:1048:60  */
  assign n4148_o = ~dp_write_stream_rrrrr;
  /* ../../HW/src/pcore/core.vhd:1048:34  */
  assign n4149_o = n4148_o ? dp_writedata_rrrrr : stream_write_output;
  /* ../../HW/src/pcore/core.vhd:1090:32  */
  assign gen_cell_n1_cell_i_n4152 = gen_cell_n1_cell_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1091:33  */
  assign gen_cell_n1_cell_i_n4153 = gen_cell_n1_cell_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1092:35  */
  assign gen_cell_n1_cell_i_n4154 = gen_cell_n1_cell_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1093:34  */
  assign gen_cell_n1_cell_i_n4155 = gen_cell_n1_cell_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1094:38  */
  assign gen_cell_n1_cell_i_n4156 = gen_cell_n1_cell_i_dp_readdata_valid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1095:38  */
  assign gen_cell_n1_cell_i_n4157 = gen_cell_n1_cell_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1096:37  */
  assign gen_cell_n1_cell_i_n4158 = gen_cell_n1_cell_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1098:33  */
  assign gen_cell_n1_cell_i_n4160 = gen_cell_n1_cell_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1099:36  */
  assign gen_cell_n1_cell_i_n4161 = gen_cell_n1_cell_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1110:32  */
  assign n4162_o = enable[3:0];
  /* ../../HW/src/pcore/core.vhd:1120:29  */
  assign gen_cell_n1_cell_i_n4163 = gen_cell_n1_cell_i_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1121:29  */
  assign gen_cell_n1_cell_i_n4164 = gen_cell_n1_cell_i_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  cell_0 gen_cell_n1_cell_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .dp_rd_vm_in(dp_rd_vm_r),
    .dp_wr_vm_in(dp_wr_vm_rrrrr),
    .dp_code_in(dp_code_rrrrr),
    .dp_rd_addr_in(dp_rd_addr_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_r),
    .dp_rd_fork_in(n4150_o),
    .dp_rd_share_in(dp_rd_share_r),
    .dp_wr_addr_in(dp_wr_addr_rrrrr),
    .dp_wr_addr_step_in(dp_wr_addr_step_rrrrr),
    .dp_wr_fork_in(n4151_o),
    .dp_wr_share_in(dp_wr_share_rrrrr),
    .dp_wr_mcast_in(dp_wr_mcast_rrrrr),
    .dp_write_in(dp_write_rrrrr),
    .dp_write_gen_valid_in(dp_write_gen_valid_rrrrr),
    .dp_write_vector_in(dp_write_vector_rrrrr),
    .dp_write_scatter_in(dp_write_scatter_rrrrr),
    .dp_read_in(dp_read_r),
    .dp_read_vector_in(dp_read_vector_r),
    .dp_read_scatter_in(dp_read_scatter_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_r),
    .dp_read_data_flow_in(dp_read_data_flow_r),
    .dp_read_data_type_in(dp_read_data_type_r),
    .dp_read_stream_in(dp_read_stream_r),
    .dp_read_stream_id_in(dp_read_stream_id_r),
    .dp_writedata_in(writedata2),
    .dp_config_in(dp_config_rrrrr),
    .instruction_mu_in(instruction_mu),
    .instruction_imu_in(instruction_imu),
    .instruction_mu_valid_in(instruction_mu_valid),
    .instruction_imu_valid_in(instruction_imu_valid),
    .vm_in(vm),
    .data_model_in(data_model),
    .enable_in(n4162_o),
    .tid_in(tid),
    .tid_valid1_in(tid_valid1),
    .pre_tid_in(pre_tid),
    .pre_tid_valid1_in(pre_tid_valid1),
    .pre_pre_tid_in(pre_pre_tid),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1),
    .pre_pre_vm_in(pre_pre_vm),
    .pre_pre_data_model_in(pre_pre_data_model),
    .pre_iregister_auto_in(pre_iregister_auto),
    .dp_readdata_out(gen_cell_n1_cell_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_cell_n1_cell_i_dp_readdata_vm_out),
    .dp_read_vector_out(gen_cell_n1_cell_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_cell_n1_cell_i_dp_read_vaddr_out),
    .dp_readdata_valid_out(gen_cell_n1_cell_i_dp_readdata_valid_out),
    .dp_read_gen_valid_out(gen_cell_n1_cell_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_cell_n1_cell_i_dp_read_data_flow_out),
    .dp_read_data_type_out(),
    .dp_read_stream_out(gen_cell_n1_cell_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_cell_n1_cell_i_dp_read_stream_id_out),
    .i_y_neg_out(gen_cell_n1_cell_i_i_y_neg_out),
    .i_y_zero_out(gen_cell_n1_cell_i_i_y_zero_out));
  /* ../../HW/src/pcore/core.vhd:1090:32  */
  assign gen_cell_n2_cell_i_n4191 = gen_cell_n2_cell_i_dp_readdata_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1091:33  */
  assign gen_cell_n2_cell_i_n4192 = gen_cell_n2_cell_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1092:35  */
  assign gen_cell_n2_cell_i_n4193 = gen_cell_n2_cell_i_dp_read_vector_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1093:34  */
  assign gen_cell_n2_cell_i_n4194 = gen_cell_n2_cell_i_dp_read_vaddr_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1094:38  */
  assign gen_cell_n2_cell_i_n4195 = gen_cell_n2_cell_i_dp_readdata_valid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1095:38  */
  assign gen_cell_n2_cell_i_n4196 = gen_cell_n2_cell_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1096:37  */
  assign gen_cell_n2_cell_i_n4197 = gen_cell_n2_cell_i_dp_read_data_flow_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1098:33  */
  assign gen_cell_n2_cell_i_n4199 = gen_cell_n2_cell_i_dp_read_stream_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1099:36  */
  assign gen_cell_n2_cell_i_n4200 = gen_cell_n2_cell_i_dp_read_stream_id_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1110:32  */
  assign n4201_o = enable[7:4];
  /* ../../HW/src/pcore/core.vhd:1120:29  */
  assign gen_cell_n2_cell_i_n4202 = gen_cell_n2_cell_i_i_y_neg_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1121:29  */
  assign gen_cell_n2_cell_i_n4203 = gen_cell_n2_cell_i_i_y_zero_out; // (signal)
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  cell_1 gen_cell_n2_cell_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .dp_rd_vm_in(dp_rd_vm_r),
    .dp_wr_vm_in(dp_wr_vm_rrrrr),
    .dp_code_in(dp_code_rrrrr),
    .dp_rd_addr_in(dp_rd_addr_r),
    .dp_rd_addr_step_in(dp_rd_addr_step_r),
    .dp_rd_fork_in(n4189_o),
    .dp_rd_share_in(dp_rd_share_r),
    .dp_wr_addr_in(dp_wr_addr_rrrrr),
    .dp_wr_addr_step_in(dp_wr_addr_step_rrrrr),
    .dp_wr_fork_in(n4190_o),
    .dp_wr_share_in(dp_wr_share_rrrrr),
    .dp_wr_mcast_in(dp_wr_mcast_rrrrr),
    .dp_write_in(dp_write_rrrrr),
    .dp_write_gen_valid_in(dp_write_gen_valid_rrrrr),
    .dp_write_vector_in(dp_write_vector_rrrrr),
    .dp_write_scatter_in(dp_write_scatter_rrrrr),
    .dp_read_in(dp_read_r),
    .dp_read_vector_in(dp_read_vector_r),
    .dp_read_scatter_in(dp_read_scatter_r),
    .dp_read_gen_valid_in(dp_read_gen_valid_r),
    .dp_read_data_flow_in(dp_read_data_flow_r),
    .dp_read_data_type_in(dp_read_data_type_r),
    .dp_read_stream_in(dp_read_stream_r),
    .dp_read_stream_id_in(dp_read_stream_id_r),
    .dp_writedata_in(writedata2),
    .dp_config_in(dp_config_rrrrr),
    .instruction_mu_in(instruction_mu),
    .instruction_imu_in(instruction_imu),
    .instruction_mu_valid_in(instruction_mu_valid),
    .instruction_imu_valid_in(instruction_imu_valid),
    .vm_in(vm),
    .data_model_in(data_model),
    .enable_in(n4201_o),
    .tid_in(tid),
    .tid_valid1_in(tid_valid1),
    .pre_tid_in(pre_tid),
    .pre_tid_valid1_in(pre_tid_valid1),
    .pre_pre_tid_in(pre_pre_tid),
    .pre_pre_tid_valid1_in(pre_pre_tid_valid1),
    .pre_pre_vm_in(pre_pre_vm),
    .pre_pre_data_model_in(pre_pre_data_model),
    .pre_iregister_auto_in(pre_iregister_auto),
    .dp_readdata_out(gen_cell_n2_cell_i_dp_readdata_out),
    .dp_readdata_vm_out(gen_cell_n2_cell_i_dp_readdata_vm_out),
    .dp_read_vector_out(gen_cell_n2_cell_i_dp_read_vector_out),
    .dp_read_vaddr_out(gen_cell_n2_cell_i_dp_read_vaddr_out),
    .dp_readdata_valid_out(gen_cell_n2_cell_i_dp_readdata_valid_out),
    .dp_read_gen_valid_out(gen_cell_n2_cell_i_dp_read_gen_valid_out),
    .dp_read_data_flow_out(gen_cell_n2_cell_i_dp_read_data_flow_out),
    .dp_read_data_type_out(),
    .dp_read_stream_out(gen_cell_n2_cell_i_dp_read_stream_out),
    .dp_read_stream_id_out(gen_cell_n2_cell_i_dp_read_stream_id_out),
    .i_y_neg_out(gen_cell_n2_cell_i_i_y_neg_out),
    .i_y_zero_out(gen_cell_n2_cell_i_i_y_zero_out));
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4228_q <= 3'b000;
    else
      n4228_q <= n3676_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4229_q <= 3'b000;
    else
      n4229_q <= dp_write_vector_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4230_q <= 3'b000;
    else
      n4230_q <= dp_write_vector_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4231_q <= 3'b000;
    else
      n4231_q <= dp_write_vector_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4232_q <= 3'b000;
    else
      n4232_q <= dp_write_vector_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4233_q <= 2'b00;
    else
      n4233_q <= n3678_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4234_q <= 2'b00;
    else
      n4234_q <= dp_write_scatter_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4235_q <= 2'b00;
    else
      n4235_q <= dp_write_scatter_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4236_q <= 2'b00;
    else
      n4236_q <= dp_write_scatter_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4237_q <= 2'b00;
    else
      n4237_q <= dp_write_scatter_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4238_q <= 1'b0;
    else
      n4238_q <= n3680_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4239_q <= 1'b0;
    else
      n4239_q <= dp_wr_vm_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4240_q <= 1'b0;
    else
      n4240_q <= dp_wr_vm_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4241_q <= 1'b0;
    else
      n4241_q <= dp_wr_vm_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4242_q <= 1'b0;
    else
      n4242_q <= dp_wr_vm_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4243_q <= 1'b0;
    else
      n4243_q <= n3682_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4244_q <= 1'b0;
    else
      n4244_q <= dp_code_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4245_q <= 1'b0;
    else
      n4245_q <= dp_code_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4246_q <= 1'b0;
    else
      n4246_q <= dp_code_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4247_q <= 1'b0;
    else
      n4247_q <= dp_code_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4248_q <= 1'b0;
    else
      n4248_q <= n3685_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4249_q <= 1'b0;
    else
      n4249_q <= dp_config_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4250_q <= 1'b0;
    else
      n4250_q <= dp_config_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4251_q <= 1'b0;
    else
      n4251_q <= dp_config_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4252_q <= 1'b0;
    else
      n4252_q <= dp_config_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4253_q <= 22'b0000000000000000000000;
    else
      n4253_q <= n3734_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4254_q <= 22'b0000000000000000000000;
    else
      n4254_q <= dp_wr_addr_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4255_q <= 22'b0000000000000000000000;
    else
      n4255_q <= dp_wr_addr_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4256_q <= 22'b0000000000000000000000;
    else
      n4256_q <= dp_wr_addr_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4257_q <= 22'b0000000000000000000000;
    else
      n4257_q <= dp_wr_addr_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4258_q <= 22'b0000000000000000000000;
    else
      n4258_q <= n3691_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4259_q <= 22'b0000000000000000000000;
    else
      n4259_q <= dp_wr_addr_step_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4260_q <= 22'b0000000000000000000000;
    else
      n4260_q <= dp_wr_addr_step_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4261_q <= 22'b0000000000000000000000;
    else
      n4261_q <= dp_wr_addr_step_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4262_q <= 22'b0000000000000000000000;
    else
      n4262_q <= dp_wr_addr_step_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4263_q <= 1'b0;
    else
      n4263_q <= n3693_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4264_q <= 1'b0;
    else
      n4264_q <= dp_wr_share_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4265_q <= 1'b0;
    else
      n4265_q <= dp_wr_share_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4266_q <= 1'b0;
    else
      n4266_q <= dp_wr_share_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4267_q <= 1'b0;
    else
      n4267_q <= dp_wr_share_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4268_q <= 1'b0;
    else
      n4268_q <= n3695_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4269_q <= 1'b0;
    else
      n4269_q <= dp_write_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4270_q <= 1'b0;
    else
      n4270_q <= dp_write_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4271_q <= 1'b0;
    else
      n4271_q <= dp_write_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4272_q <= 1'b0;
    else
      n4272_q <= dp_write_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4273_q <= 1'b0;
    else
      n4273_q <= n3697_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4274_q <= 1'b0;
    else
      n4274_q <= dp_write_gen_valid_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4275_q <= 1'b0;
    else
      n4275_q <= dp_write_gen_valid_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4276_q <= 1'b0;
    else
      n4276_q <= dp_write_gen_valid_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4277_q <= 1'b0;
    else
      n4277_q <= dp_write_gen_valid_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4278_q <= 6'b111111;
    else
      n4278_q <= n3699_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4279_q <= 6'b111111;
    else
      n4279_q <= dp_wr_mcast_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4280_q <= 6'b111111;
    else
      n4280_q <= dp_wr_mcast_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4281_q <= 6'b111111;
    else
      n4281_q <= dp_wr_mcast_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4282_q <= 6'b111111;
    else
      n4282_q <= dp_wr_mcast_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4283_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4283_q <= n3702_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4284_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4284_q <= dp_writedata_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4285_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4285_q <= dp_writedata_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4286_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4286_q <= dp_writedata_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4287_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4287_q <= dp_writedata_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  assign n4288_o = n3597_o ? n3599_o : dp_stream_read_req_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4289_q <= 8'b00000000;
    else
      n4289_q <= n4288_o;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  assign n4290_o = dp_read_stream2_r ? n3261_o : dp_stream_read_done_r;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4291_q <= 8'b00000000;
    else
      n4291_q <= n4290_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4292_q <= 3'b000;
    else
      n4292_q <= dp_read_vector_in;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4293_q <= 2'b00;
    else
      n4293_q <= dp_read_scatter_in;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4294_q <= 2'b00;
    else
      n4294_q <= dp_read_data_flow_in;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4295_q <= 2'b00;
    else
      n4295_q <= dp_read_data_flow;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4296_q <= 2'b00;
    else
      n4296_q <= dp_read_data_flow2_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4297_q <= 2'b00;
    else
      n4297_q <= dp_read_data_flow2_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4298_q <= 2'b00;
    else
      n4298_q <= dp_read_data_flow2_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4299_q <= 2'b00;
    else
      n4299_q <= dp_read_data_flow2_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4300_q <= 2'b00;
    else
      n4300_q <= dp_read_data_type_in;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4306_q <= 1'b0;
    else
      n4306_q <= dp_read_stream_in;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4307_q <= 2'b00;
    else
      n4307_q <= dp_read_stream_id_in;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4308_q <= 2'b00;
    else
      n4308_q <= dp_read_stream_id;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4309_q <= 1'b0;
    else
      n4309_q <= dp_rd_vm;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4310_q <= 2'b00;
    else
      n4310_q <= busy;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4311_q <= 1'b0;
    else
      n4311_q <= ready;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4313_q <= 22'b0000000000000000000000;
    else
      n4313_q <= dp_rd_addr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4314_q <= 22'b0000000000000000000000;
    else
      n4314_q <= dp_rd_addr_step;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4315_q <= 1'b0;
    else
      n4315_q <= dp_rd_share;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4316_q <= 1'b0;
    else
      n4316_q <= dp_core_read;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4317_q <= 1'b0;
    else
      n4317_q <= dp_read_gen_valid_in;
  /* ../../HW/src/pcore/core.vhd:617:5  */
  assign n4318_o = {gen_cell_n2_cell_i_n4195, gen_cell_n1_cell_i_n4156};
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4319_o = gen_cell_n1_cell_i_n4157;
  assign n4319_o = gen_cell_n2_cell_i_n4196;
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4320_o = gen_cell_n1_cell_i_n4153;
  assign n4320_o = gen_cell_n2_cell_i_n4192;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4321_q <= 1'b0;
    else
      n4321_q <= dp_readdata_vm;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4322_q <= 1'b0;
    else
      n4322_q <= dp_readdata_vm_r;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4323_q <= 1'b0;
    else
      n4323_q <= dp_readdata_vm_rr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4324_q <= 1'b0;
    else
      n4324_q <= dp_readdata_vm_rrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4325_q <= 1'b0;
    else
      n4325_q <= dp_readdata_vm_rrrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4326_q <= 1'b0;
    else
      n4326_q <= dp_readdata_vm_rrrrr;
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4327_o = gen_cell_n1_cell_i_n4158;
  assign n4327_o = gen_cell_n2_cell_i_n4197;
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4329_o = gen_cell_n1_cell_i_n4160;
  assign n4329_o = gen_cell_n2_cell_i_n4199;
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4330_o = gen_cell_n1_cell_i_n4161;
  assign n4330_o = gen_cell_n2_cell_i_n4200;
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4331_o = gen_cell_n1_cell_i_n4152;
  assign n4331_o = gen_cell_n2_cell_i_n4191;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4332_q <= 1'b0;
    else
      n4332_q <= dp_readdatavalid;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4333_q <= 1'b0;
    else
      n4333_q <= dp_readdatavalid2_r;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4334_q <= 1'b0;
    else
      n4334_q <= dp_readdatavalid2_rr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4335_q <= 1'b0;
    else
      n4335_q <= dp_readdatavalid2_rrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4336_q <= 1'b0;
    else
      n4336_q <= dp_readdatavalid2_rrrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4337_q <= 1'b0;
    else
      n4337_q <= dp_readdatavalid2_rrrrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4338_q <= 1'b0;
    else
      n4338_q <= dp_read_gen_valid;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4339_q <= 1'b0;
    else
      n4339_q <= dp_read_gen_valid2_r;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4340_q <= 1'b0;
    else
      n4340_q <= dp_read_gen_valid2_rr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4341_q <= 1'b0;
    else
      n4341_q <= dp_read_gen_valid2_rrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4342_q <= 1'b0;
    else
      n4342_q <= dp_read_gen_valid2_rrrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4343_q <= 1'b0;
    else
      n4343_q <= dp_read_gen_valid2_rrrrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4344_q <= 1'b0;
    else
      n4344_q <= n3259_o;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4345_q <= 1'b0;
    else
      n4345_q <= dp_read_stream2_r;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4346_q <= 1'b0;
    else
      n4346_q <= dp_read_stream2_rr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4347_q <= 1'b0;
    else
      n4347_q <= dp_read_stream2_rrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4348_q <= 1'b0;
    else
      n4348_q <= dp_read_stream2_rrrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4350_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4350_q <= dp_readdata2;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4351_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4351_q <= dp_readdata2_r;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4352_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4352_q <= dp_readdata2_rr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4353_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4353_q <= dp_readdata2_rrr;
  /* ../../HW/src/pcore/core.vhd:531:8  */
  always @(posedge clock_in or posedge n3255_o)
    if (n3255_o)
      n4354_q <= 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n4354_q <= dp_readdata2_rrrr;
  /* ../../HW/src/pcore/core.vhd:492:5  */
  assign n4356_o = {gen_stream_n8_stream_i_n3069, gen_stream_n7_stream_i_n3065, gen_stream_n6_stream_i_n3061, gen_stream_n5_stream_i_n3057, gen_stream_n4_stream_i_n3053, gen_stream_n3_stream_i_n3049, gen_stream_n2_stream_i_n3045, gen_stream_n1_stream_i_n3041};
  /* ../../HW/src/pcore/core.vhd:492:5  */
  assign n4357_o = {gen_stream_1_n8_stream_i1_n3101, gen_stream_1_n7_stream_i1_n3097, gen_stream_1_n6_stream_i1_n3093, gen_stream_1_n5_stream_i1_n3089, gen_stream_1_n4_stream_i1_n3085, gen_stream_1_n3_stream_i1_n3081, gen_stream_1_n2_stream_i1_n3077, gen_stream_1_n1_stream_i1_n3073};
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4358_o = gen_cell_n1_cell_i_n4154;
  assign n4358_o = gen_cell_n2_cell_i_n4193;
  /* ../../HW/src/pcore/core.vhd:1056:1  */
  assign n4359_o = gen_cell_n1_cell_i_n4155;
  assign n4359_o = gen_cell_n2_cell_i_n4194;
  /* ../../HW/src/pcore/core.vhd:448:9  */
  always @(posedge clock_in or posedge n3130_o)
    if (n3130_o)
      n4360_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n4360_q <= n3216_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4361_q <= 1'b0;
    else
      n4361_q <= 1'b0;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4362_q <= 1'b0;
    else
      n4362_q <= 1'b0;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4363_q <= 1'b0;
    else
      n4363_q <= n3704_o;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4364_q <= 1'b0;
    else
      n4364_q <= dp_write_stream_r;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4365_q <= 1'b0;
    else
      n4365_q <= dp_write_stream_rr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4366_q <= 1'b0;
    else
      n4366_q <= dp_write_stream_rrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4367_q <= 1'b0;
    else
      n4367_q <= dp_write_stream_rrrr;
  /* ../../HW/src/pcore/core.vhd:727:9  */
  always @(posedge clock_in or posedge n3595_o)
    if (n3595_o)
      n4368_q <= 2'b00;
    else
      n4368_q <= n3706_o;
  /* ../../HW/src/pcore/core.vhd:617:5  */
  assign n4369_o = {gen_cell_n2_cell_i_n4202, gen_cell_n1_cell_i_n4163};
  /* ../../HW/src/pcore/core.vhd:617:5  */
  assign n4370_o = {gen_cell_n2_cell_i_n4203, gen_cell_n1_cell_i_n4164};
endmodule

module dp_core
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  [11:0] bus_waddr_in,
   input  [11:0] bus_raddr_in,
   input  bus_write_in,
   input  bus_read_in,
   input  [31:0] bus_writedata_in,
   input  readmaster1_readdatavalid_in,
   input  readmaster1_readdatavalid_vm_in,
   input  [63:0] readmaster1_readdata_in,
   input  readmaster1_wait_request_in,
   input  writemaster1_wait_request_in,
   input  [47:0] writemaster1_counter_in,
   input  readmaster2_readdatavalid_in,
   input  readmaster2_readdatavalid_vm_in,
   input  [63:0] readmaster2_readdata_in,
   input  readmaster2_wait_request_in,
   input  writemaster2_wait_request_in,
   input  [47:0] writemaster2_counter_in,
   input  readmaster3_readdatavalid_in,
   input  readmaster3_readdatavalid_vm_in,
   input  [63:0] readmaster3_readdata_in,
   input  readmaster3_wait_request_in,
   input  writemaster3_wait_request_in,
   input  [23:0] writemaster3_counter_in,
   input  [1:0] task_busy_in,
   input  task_ready_in,
   input  [71:0] bar_in,
   input  ddr_tx_busy_in,
   output [31:0] bus_readdata_out,
   output bus_readdatavalid_out,
   output bus_writewait_out,
   output bus_readwait_out,
   output [21:0] readmaster1_addr_out,
   output readmaster1_fork_out,
   output readmaster1_addr_mode_out,
   output readmaster1_cs_out,
   output readmaster1_read_out,
   output readmaster1_read_vm_out,
   output [1:0] readmaster1_read_data_flow_out,
   output readmaster1_read_stream_out,
   output [1:0] readmaster1_read_stream_id_out,
   output [2:0] readmaster1_read_vector_out,
   output [1:0] readmaster1_read_scatter_out,
   output [4:0] readmaster1_burstlen_out,
   output [1:0] readmaster1_bus_id_out,
   output [1:0] readmaster1_data_type_out,
   output [1:0] readmaster1_data_model_out,
   output [21:0] writemaster1_addr_out,
   output writemaster1_fork_out,
   output writemaster1_addr_mode_out,
   output writemaster1_vm_out,
   output [5:0] writemaster1_mcast_out,
   output writemaster1_cs_out,
   output writemaster1_write_out,
   output [1:0] writemaster1_write_data_flow_out,
   output [2:0] writemaster1_write_vector_out,
   output writemaster1_write_stream_out,
   output [1:0] writemaster1_write_stream_id_out,
   output [1:0] writemaster1_write_scatter_out,
   output [63:0] writemaster1_writedata_out,
   output [4:0] writemaster1_burstlen_out,
   output [1:0] writemaster1_bus_id_out,
   output [1:0] writemaster1_data_type_out,
   output [1:0] writemaster1_data_model_out,
   output writemaster1_thread_out,
   output [17:0] readmaster2_addr_out,
   output readmaster2_fork_out,
   output readmaster2_cs_out,
   output readmaster2_read_out,
   output readmaster2_read_vm_out,
   output [2:0] readmaster2_read_vector_out,
   output [1:0] readmaster2_read_scatter_out,
   output [4:0] readmaster2_burstlen_out,
   output [1:0] readmaster2_bus_id_out,
   output [17:0] writemaster2_addr_out,
   output writemaster2_fork_out,
   output writemaster2_cs_out,
   output writemaster2_write_out,
   output writemaster2_vm_out,
   output [2:0] writemaster2_write_vector_out,
   output [1:0] writemaster2_write_scatter_out,
   output [63:0] writemaster2_writedata_out,
   output [4:0] writemaster2_burstlen_out,
   output [1:0] writemaster2_bus_id_out,
   output writemaster2_thread_out,
   output [31:0] readmaster3_addr_out,
   output readmaster3_cs_out,
   output readmaster3_read_out,
   output readmaster3_read_vm_out,
   output [2:0] readmaster3_read_vector_out,
   output [1:0] readmaster3_read_scatter_out,
   output [3:0] readmaster3_read_start_out,
   output [3:0] readmaster3_read_end_out,
   output [4:0] readmaster3_burstlen_out,
   output [1:0] readmaster3_bus_id_out,
   output [15:0] readmaster3_filler_data_out,
   output [31:0] writemaster3_addr_out,
   output writemaster3_cs_out,
   output writemaster3_write_out,
   output writemaster3_vm_out,
   output [2:0] writemaster3_write_vector_out,
   output [1:0] writemaster3_write_scatter_out,
   output [3:0] writemaster3_write_end_out,
   output [63:0] writemaster3_writedata_out,
   output [4:0] writemaster3_burstlen_out,
   output [8:0] writemaster3_burstlen2_out,
   output [4:0] writemaster3_burstlen3_out,
   output [1:0] writemaster3_bus_id_out,
   output writemaster3_thread_out,
   output [15:0] writemaster3_filler_data_out,
   output [10:0] task_start_addr_out,
   output task_out,
   output task_vm_out,
   output [4:0] task_pcore_out,
   output task_lockstep_out,
   output [3:0] task_tid_mask_out,
   output [27:0] task_iregister_auto_out,
   output [1:0] task_data_model_out,
   output [1:0] task_busy_out,
   output indication_avail_out);
  wire [1:0] task_busy;
  wire task_ready;
  wire \task ;
  wire [4:0] task_pcore;
  wire task_lockstep;
  wire [3:0] task_tid_mask;
  wire [27:0] task_iregister_auto;
  wire [1:0] task_data_model;
  wire [10:0] task_start_addr;
  wire task_vm;
  reg [4:0] task_pcore_r;
  wire task_lockstep_r;
  wire [3:0] task_tid_mask_r;
  wire [27:0] task_iregister_auto_r;
  wire [1:0] task_data_model_r;
  wire [10:0] task_start_addr_r;
  wire task_r;
  wire task_rr;
  wire task_rrr;
  wire task_rrrr;
  wire task_rrrrr;
  wire task_rrrrrr;
  wire task_rrrrrrr;
  wire task_rrrrrrrr;
  wire task_vm_r;
  wire task_vm_rr;
  wire task_vm_rrr;
  wire task_vm_rrrr;
  wire task_vm_rrrrr;
  wire task_vm_rrrrrr;
  wire task_vm_rrrrrrr;
  wire task_vm_rrrrrrrr;
  wire task_busy_r;
  wire task_1_busy_r;
  wire task_0_busy_r;
  wire [31:0] dp0_i_n2576;
  wire dp0_i_n2577;
  wire dp0_i_n2578;
  wire dp0_i_n2579;
  wire [21:0] dp0_i_n2580;
  wire dp0_i_n2581;
  wire dp0_i_n2582;
  wire dp0_i_n2583;
  wire dp0_i_n2584;
  wire dp0_i_n2585;
  wire [1:0] dp0_i_n2586;
  wire dp0_i_n2587;
  wire [1:0] dp0_i_n2588;
  wire [2:0] dp0_i_n2589;
  wire [1:0] dp0_i_n2590;
  wire [4:0] dp0_i_n2591;
  wire [1:0] dp0_i_n2592;
  wire [1:0] dp0_i_n2593;
  wire [1:0] dp0_i_n2594;
  wire [21:0] dp0_i_n2595;
  wire dp0_i_n2596;
  wire dp0_i_n2597;
  wire dp0_i_n2598;
  wire [5:0] dp0_i_n2599;
  wire dp0_i_n2600;
  wire dp0_i_n2601;
  wire [1:0] dp0_i_n2602;
  wire [2:0] dp0_i_n2603;
  wire dp0_i_n2604;
  wire [1:0] dp0_i_n2605;
  wire [1:0] dp0_i_n2606;
  wire [63:0] dp0_i_n2607;
  wire [4:0] dp0_i_n2608;
  wire [1:0] dp0_i_n2609;
  wire [1:0] dp0_i_n2610;
  wire [1:0] dp0_i_n2611;
  wire dp0_i_n2612;
  wire [17:0] dp0_i_n2613;
  wire dp0_i_n2614;
  wire dp0_i_n2615;
  wire dp0_i_n2616;
  wire dp0_i_n2617;
  wire [2:0] dp0_i_n2618;
  wire [1:0] dp0_i_n2619;
  wire [4:0] dp0_i_n2620;
  wire [1:0] dp0_i_n2621;
  wire [17:0] dp0_i_n2622;
  wire dp0_i_n2623;
  wire dp0_i_n2624;
  wire dp0_i_n2625;
  wire dp0_i_n2626;
  wire [2:0] dp0_i_n2627;
  wire [1:0] dp0_i_n2628;
  wire [63:0] dp0_i_n2629;
  wire [4:0] dp0_i_n2630;
  wire [1:0] dp0_i_n2631;
  wire dp0_i_n2632;
  wire [31:0] dp0_i_n2633;
  wire dp0_i_n2634;
  wire dp0_i_n2635;
  wire dp0_i_n2636;
  wire [2:0] dp0_i_n2637;
  wire [1:0] dp0_i_n2638;
  wire [3:0] dp0_i_n2639;
  wire [3:0] dp0_i_n2640;
  wire [4:0] dp0_i_n2641;
  wire [1:0] dp0_i_n2642;
  wire [15:0] dp0_i_n2643;
  wire [31:0] dp0_i_n2644;
  wire dp0_i_n2645;
  wire dp0_i_n2646;
  wire dp0_i_n2647;
  wire [2:0] dp0_i_n2648;
  wire [1:0] dp0_i_n2649;
  wire [3:0] dp0_i_n2650;
  wire [63:0] dp0_i_n2651;
  wire [4:0] dp0_i_n2652;
  wire [8:0] dp0_i_n2653;
  wire [4:0] dp0_i_n2654;
  wire [1:0] dp0_i_n2655;
  wire dp0_i_n2656;
  wire [10:0] dp0_i_n2657;
  wire dp0_i_n2658;
  wire dp0_i_n2660;
  wire [4:0] dp0_i_n2661;
  wire dp0_i_n2662;
  wire [3:0] dp0_i_n2663;
  wire [27:0] dp0_i_n2664;
  wire [1:0] dp0_i_n2665;
  wire dp0_i_n2666;
  wire [31:0] dp0_i_bus_readdata_out;
  wire dp0_i_bus_readdatavalid_out;
  wire dp0_i_bus_writewait_out;
  wire dp0_i_bus_readwait_out;
  wire [21:0] dp0_i_readmaster1_addr_out;
  wire dp0_i_readmaster1_fork_out;
  wire dp0_i_readmaster1_addr_mode_out;
  wire dp0_i_readmaster1_cs_out;
  wire dp0_i_readmaster1_read_out;
  wire dp0_i_readmaster1_read_vm_out;
  wire [1:0] dp0_i_readmaster1_read_data_flow_out;
  wire dp0_i_readmaster1_read_stream_out;
  wire [1:0] dp0_i_readmaster1_read_stream_id_out;
  wire [2:0] dp0_i_readmaster1_read_vector_out;
  wire [1:0] dp0_i_readmaster1_read_scatter_out;
  wire [4:0] dp0_i_readmaster1_burstlen_out;
  wire [1:0] dp0_i_readmaster1_bus_id_out;
  wire [1:0] dp0_i_readmaster1_data_type_out;
  wire [1:0] dp0_i_readmaster1_data_model_out;
  wire [21:0] dp0_i_writemaster1_addr_out;
  wire dp0_i_writemaster1_fork_out;
  wire dp0_i_writemaster1_addr_mode_out;
  wire dp0_i_writemaster1_vm_out;
  wire [5:0] dp0_i_writemaster1_mcast_out;
  wire dp0_i_writemaster1_cs_out;
  wire dp0_i_writemaster1_write_out;
  wire [1:0] dp0_i_writemaster1_write_data_flow_out;
  wire [2:0] dp0_i_writemaster1_write_vector_out;
  wire dp0_i_writemaster1_write_stream_out;
  wire [1:0] dp0_i_writemaster1_write_stream_id_out;
  wire [1:0] dp0_i_writemaster1_write_scatter_out;
  wire [63:0] dp0_i_writemaster1_writedata_out;
  wire [4:0] dp0_i_writemaster1_burstlen_out;
  wire [1:0] dp0_i_writemaster1_bus_id_out;
  wire [1:0] dp0_i_writemaster1_data_type_out;
  wire [1:0] dp0_i_writemaster1_data_model_out;
  wire dp0_i_writemaster1_thread_out;
  wire [17:0] dp0_i_readmaster2_addr_out;
  wire dp0_i_readmaster2_fork_out;
  wire dp0_i_readmaster2_cs_out;
  wire dp0_i_readmaster2_read_out;
  wire dp0_i_readmaster2_read_vm_out;
  wire [2:0] dp0_i_readmaster2_read_vector_out;
  wire [1:0] dp0_i_readmaster2_read_scatter_out;
  wire [4:0] dp0_i_readmaster2_burstlen_out;
  wire [1:0] dp0_i_readmaster2_bus_id_out;
  wire [17:0] dp0_i_writemaster2_addr_out;
  wire dp0_i_writemaster2_vm_out;
  wire dp0_i_writemaster2_fork_out;
  wire dp0_i_writemaster2_cs_out;
  wire dp0_i_writemaster2_write_out;
  wire [2:0] dp0_i_writemaster2_write_vector_out;
  wire [1:0] dp0_i_writemaster2_write_scatter_out;
  wire [63:0] dp0_i_writemaster2_writedata_out;
  wire [4:0] dp0_i_writemaster2_burstlen_out;
  wire [1:0] dp0_i_writemaster2_bus_id_out;
  wire dp0_i_writemaster2_thread_out;
  wire [31:0] dp0_i_readmaster3_addr_out;
  wire dp0_i_readmaster3_cs_out;
  wire dp0_i_readmaster3_read_out;
  wire dp0_i_readmaster3_read_vm_out;
  wire [2:0] dp0_i_readmaster3_read_vector_out;
  wire [1:0] dp0_i_readmaster3_read_scatter_out;
  wire [3:0] dp0_i_readmaster3_read_start_out;
  wire [3:0] dp0_i_readmaster3_read_end_out;
  wire [4:0] dp0_i_readmaster3_burstlen_out;
  wire [1:0] dp0_i_readmaster3_bus_id_out;
  wire [15:0] dp0_i_readmaster3_filler_data_out;
  wire [31:0] dp0_i_writemaster3_addr_out;
  wire dp0_i_writemaster3_cs_out;
  wire dp0_i_writemaster3_write_out;
  wire dp0_i_writemaster3_vm_out;
  wire [2:0] dp0_i_writemaster3_write_vector_out;
  wire [1:0] dp0_i_writemaster3_write_scatter_out;
  wire [3:0] dp0_i_writemaster3_write_end_out;
  wire [63:0] dp0_i_writemaster3_writedata_out;
  wire [4:0] dp0_i_writemaster3_burstlen_out;
  wire [8:0] dp0_i_writemaster3_burstlen2_out;
  wire [4:0] dp0_i_writemaster3_burstlen3_out;
  wire [1:0] dp0_i_writemaster3_bus_id_out;
  wire dp0_i_writemaster3_thread_out;
  wire [10:0] dp0_i_task_start_addr_out;
  wire dp0_i_task_out;
  wire dp0_i_task_pending_out;
  wire dp0_i_task_vm_out;
  wire [4:0] dp0_i_task_pcore_out;
  wire dp0_i_task_lockstep_out;
  wire [3:0] dp0_i_task_tid_mask_out;
  wire [27:0] dp0_i_task_iregister_auto_out;
  wire [1:0] dp0_i_task_data_model_out;
  wire dp0_i_indication_avail_out;
  wire n2850_o;
  wire n2851_o;
  wire n2852_o;
  wire n2855_o;
  wire n2856_o;
  wire n2857_o;
  wire n2860_o;
  wire n2861_o;
  wire n2862_o;
  wire n2866_o;
  wire n2868_o;
  wire n2869_o;
  wire n2870_o;
  wire n2871_o;
  wire n2872_o;
  wire n2873_o;
  wire n2874_o;
  wire n2875_o;
  wire n2876_o;
  wire n2877_o;
  wire n2878_o;
  wire n2879_o;
  wire n2880_o;
  wire n2881_o;
  wire n2882_o;
  wire n2883_o;
  wire n2884_o;
  wire n2885_o;
  wire n2886_o;
  wire n2887_o;
  wire n2888_o;
  wire n2889_o;
  wire n2890_o;
  wire n2891_o;
  wire n2892_o;
  wire n2893_o;
  wire n2894_o;
  wire n2895_o;
  wire n2896_o;
  wire n2897_o;
  wire n2898_o;
  wire n2899_o;
  wire n2900_o;
  wire n2901_o;
  wire n2902_o;
  wire n2903_o;
  wire n2904_o;
  wire n2905_o;
  wire n2906_o;
  wire n2907_o;
  wire n2908_o;
  wire n2909_o;
  wire n2910_o;
  wire n2911_o;
  wire n2912_o;
  wire n2913_o;
  wire n2914_o;
  wire n2915_o;
  wire n2916_o;
  wire n2917_o;
  wire n2918_o;
  wire [1:0] n2995_o;
  reg [4:0] n2996_q;
  reg n2997_q;
  reg [3:0] n2998_q;
  reg [27:0] n2999_q;
  reg [1:0] n3000_q;
  reg [10:0] n3001_q;
  reg n3002_q;
  reg n3003_q;
  reg n3004_q;
  reg n3005_q;
  reg n3006_q;
  reg n3007_q;
  reg n3008_q;
  reg n3009_q;
  reg n3010_q;
  reg n3011_q;
  reg n3012_q;
  reg n3013_q;
  reg n3014_q;
  reg n3015_q;
  reg n3016_q;
  reg n3017_q;
  reg n3018_q;
  reg n3019_q;
  reg n3020_q;
  localparam [15:0] n3021_o = 16'bZ;
  assign bus_readdata_out = dp0_i_n2576;
  assign bus_readdatavalid_out = dp0_i_n2577;
  assign bus_writewait_out = dp0_i_n2578;
  assign bus_readwait_out = dp0_i_n2579;
  assign readmaster1_addr_out = dp0_i_n2580;
  assign readmaster1_fork_out = dp0_i_n2581;
  assign readmaster1_addr_mode_out = dp0_i_n2582;
  assign readmaster1_cs_out = dp0_i_n2583;
  assign readmaster1_read_out = dp0_i_n2584;
  assign readmaster1_read_vm_out = dp0_i_n2585;
  assign readmaster1_read_data_flow_out = dp0_i_n2586;
  assign readmaster1_read_stream_out = dp0_i_n2587;
  assign readmaster1_read_stream_id_out = dp0_i_n2588;
  assign readmaster1_read_vector_out = dp0_i_n2589;
  assign readmaster1_read_scatter_out = dp0_i_n2590;
  assign readmaster1_burstlen_out = dp0_i_n2591;
  assign readmaster1_bus_id_out = dp0_i_n2592;
  assign readmaster1_data_type_out = dp0_i_n2593;
  assign readmaster1_data_model_out = dp0_i_n2594;
  assign writemaster1_addr_out = dp0_i_n2595;
  assign writemaster1_fork_out = dp0_i_n2596;
  assign writemaster1_addr_mode_out = dp0_i_n2597;
  assign writemaster1_vm_out = dp0_i_n2598;
  assign writemaster1_mcast_out = dp0_i_n2599;
  assign writemaster1_cs_out = dp0_i_n2600;
  assign writemaster1_write_out = dp0_i_n2601;
  assign writemaster1_write_data_flow_out = dp0_i_n2602;
  assign writemaster1_write_vector_out = dp0_i_n2603;
  assign writemaster1_write_stream_out = dp0_i_n2604;
  assign writemaster1_write_stream_id_out = dp0_i_n2605;
  assign writemaster1_write_scatter_out = dp0_i_n2606;
  assign writemaster1_writedata_out = dp0_i_n2607;
  assign writemaster1_burstlen_out = dp0_i_n2608;
  assign writemaster1_bus_id_out = dp0_i_n2609;
  assign writemaster1_data_type_out = dp0_i_n2610;
  assign writemaster1_data_model_out = dp0_i_n2611;
  assign writemaster1_thread_out = dp0_i_n2612;
  assign readmaster2_addr_out = dp0_i_n2613;
  assign readmaster2_fork_out = dp0_i_n2614;
  assign readmaster2_cs_out = dp0_i_n2615;
  assign readmaster2_read_out = dp0_i_n2616;
  assign readmaster2_read_vm_out = dp0_i_n2617;
  assign readmaster2_read_vector_out = dp0_i_n2618;
  assign readmaster2_read_scatter_out = dp0_i_n2619;
  assign readmaster2_burstlen_out = dp0_i_n2620;
  assign readmaster2_bus_id_out = dp0_i_n2621;
  assign writemaster2_addr_out = dp0_i_n2622;
  assign writemaster2_fork_out = dp0_i_n2623;
  assign writemaster2_cs_out = dp0_i_n2624;
  assign writemaster2_write_out = dp0_i_n2625;
  assign writemaster2_vm_out = dp0_i_n2626;
  assign writemaster2_write_vector_out = dp0_i_n2627;
  assign writemaster2_write_scatter_out = dp0_i_n2628;
  assign writemaster2_writedata_out = dp0_i_n2629;
  assign writemaster2_burstlen_out = dp0_i_n2630;
  assign writemaster2_bus_id_out = dp0_i_n2631;
  assign writemaster2_thread_out = dp0_i_n2632;
  assign readmaster3_addr_out = dp0_i_n2633;
  assign readmaster3_cs_out = dp0_i_n2634;
  assign readmaster3_read_out = dp0_i_n2635;
  assign readmaster3_read_vm_out = dp0_i_n2636;
  assign readmaster3_read_vector_out = dp0_i_n2637;
  assign readmaster3_read_scatter_out = dp0_i_n2638;
  assign readmaster3_read_start_out = dp0_i_n2639;
  assign readmaster3_read_end_out = dp0_i_n2640;
  assign readmaster3_burstlen_out = dp0_i_n2641;
  assign readmaster3_bus_id_out = dp0_i_n2642;
  assign readmaster3_filler_data_out = dp0_i_n2643;
  assign writemaster3_addr_out = dp0_i_n2644;
  assign writemaster3_cs_out = dp0_i_n2645;
  assign writemaster3_write_out = dp0_i_n2646;
  assign writemaster3_vm_out = dp0_i_n2647;
  assign writemaster3_write_vector_out = dp0_i_n2648;
  assign writemaster3_write_scatter_out = dp0_i_n2649;
  assign writemaster3_write_end_out = dp0_i_n2650;
  assign writemaster3_writedata_out = dp0_i_n2651;
  assign writemaster3_burstlen_out = dp0_i_n2652;
  assign writemaster3_burstlen2_out = dp0_i_n2653;
  assign writemaster3_burstlen3_out = dp0_i_n2654;
  assign writemaster3_bus_id_out = dp0_i_n2655;
  assign writemaster3_thread_out = dp0_i_n2656;
  assign writemaster3_filler_data_out = n3021_o;
  assign task_start_addr_out = task_start_addr_r;
  assign task_out = task_r;
  assign task_vm_out = task_vm_r;
  assign task_pcore_out = task_pcore_r;
  assign task_lockstep_out = task_lockstep_r;
  assign task_tid_mask_out = task_tid_mask_r;
  assign task_iregister_auto_out = task_iregister_auto_r;
  assign task_data_model_out = task_data_model_r;
  assign task_busy_out = task_busy;
  assign indication_avail_out = dp0_i_n2666;
  /* ../../HW/src/dp/dp_core.vhd:190:8  */
  assign task_busy = n2995_o; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:191:8  */
  assign task_ready = n2862_o; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:192:8  */
  assign \task  = dp0_i_n2658; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:194:8  */
  assign task_pcore = dp0_i_n2661; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:195:8  */
  assign task_lockstep = dp0_i_n2662; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:196:8  */
  assign task_tid_mask = dp0_i_n2663; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:197:8  */
  assign task_iregister_auto = dp0_i_n2664; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:198:8  */
  assign task_data_model = dp0_i_n2665; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:199:8  */
  assign task_start_addr = dp0_i_n2657; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:200:8  */
  assign task_vm = dp0_i_n2660; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:201:8  */
  always @*
    task_pcore_r = n2996_q; // (isignal)
  initial
    task_pcore_r = 5'b11111;
  /* ../../HW/src/dp/dp_core.vhd:202:8  */
  assign task_lockstep_r = n2997_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:203:8  */
  assign task_tid_mask_r = n2998_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:204:8  */
  assign task_iregister_auto_r = n2999_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:205:8  */
  assign task_data_model_r = n3000_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:206:8  */
  assign task_start_addr_r = n3001_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:207:8  */
  assign task_r = n3002_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:208:8  */
  assign task_rr = n3003_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:209:8  */
  assign task_rrr = n3004_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:210:8  */
  assign task_rrrr = n3005_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:211:8  */
  assign task_rrrrr = n3006_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:212:8  */
  assign task_rrrrrr = n3007_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:213:8  */
  assign task_rrrrrrr = n3008_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:214:8  */
  assign task_rrrrrrrr = n3009_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:215:8  */
  assign task_vm_r = n3010_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:216:8  */
  assign task_vm_rr = n3011_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:217:8  */
  assign task_vm_rrr = n3012_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:218:8  */
  assign task_vm_rrrr = n3013_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:219:8  */
  assign task_vm_rrrrr = n3014_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:220:8  */
  assign task_vm_rrrrrr = n3015_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:221:8  */
  assign task_vm_rrrrrrr = n3016_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:222:8  */
  assign task_vm_rrrrrrrr = n3017_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:223:8  */
  assign task_busy_r = n3018_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:224:8  */
  assign task_1_busy_r = n3019_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:225:8  */
  assign task_0_busy_r = n3020_q; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:260:27  */
  assign dp0_i_n2576 = dp0_i_bus_readdata_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:261:32  */
  assign dp0_i_n2577 = dp0_i_bus_readdatavalid_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:262:28  */
  assign dp0_i_n2578 = dp0_i_bus_writewait_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:263:27  */
  assign dp0_i_n2579 = dp0_i_bus_readwait_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:267:31  */
  assign dp0_i_n2580 = dp0_i_readmaster1_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:268:31  */
  assign dp0_i_n2581 = dp0_i_readmaster1_fork_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:269:36  */
  assign dp0_i_n2582 = dp0_i_readmaster1_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:270:29  */
  assign dp0_i_n2583 = dp0_i_readmaster1_cs_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:271:31  */
  assign dp0_i_n2584 = dp0_i_readmaster1_read_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:272:34  */
  assign dp0_i_n2585 = dp0_i_readmaster1_read_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:273:41  */
  assign dp0_i_n2586 = dp0_i_readmaster1_read_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:274:38  */
  assign dp0_i_n2587 = dp0_i_readmaster1_read_stream_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:275:41  */
  assign dp0_i_n2588 = dp0_i_readmaster1_read_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:276:38  */
  assign dp0_i_n2589 = dp0_i_readmaster1_read_vector_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:277:39  */
  assign dp0_i_n2590 = dp0_i_readmaster1_read_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:282:35  */
  assign dp0_i_n2591 = dp0_i_readmaster1_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:283:33  */
  assign dp0_i_n2592 = dp0_i_readmaster1_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:284:36  */
  assign dp0_i_n2593 = dp0_i_readmaster1_data_type_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:285:37  */
  assign dp0_i_n2594 = dp0_i_readmaster1_data_model_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:289:32  */
  assign dp0_i_n2595 = dp0_i_writemaster1_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:290:32  */
  assign dp0_i_n2596 = dp0_i_writemaster1_fork_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:291:37  */
  assign dp0_i_n2597 = dp0_i_writemaster1_addr_mode_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:292:30  */
  assign dp0_i_n2598 = dp0_i_writemaster1_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:293:33  */
  assign dp0_i_n2599 = dp0_i_writemaster1_mcast_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:294:30  */
  assign dp0_i_n2600 = dp0_i_writemaster1_cs_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:295:33  */
  assign dp0_i_n2601 = dp0_i_writemaster1_write_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:296:43  */
  assign dp0_i_n2602 = dp0_i_writemaster1_write_data_flow_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:297:40  */
  assign dp0_i_n2603 = dp0_i_writemaster1_write_vector_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:298:40  */
  assign dp0_i_n2604 = dp0_i_writemaster1_write_stream_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:299:43  */
  assign dp0_i_n2605 = dp0_i_writemaster1_write_stream_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:300:41  */
  assign dp0_i_n2606 = dp0_i_writemaster1_write_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:301:37  */
  assign dp0_i_n2607 = dp0_i_writemaster1_writedata_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:303:36  */
  assign dp0_i_n2608 = dp0_i_writemaster1_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:304:34  */
  assign dp0_i_n2609 = dp0_i_writemaster1_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:305:37  */
  assign dp0_i_n2610 = dp0_i_writemaster1_data_type_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:306:38  */
  assign dp0_i_n2611 = dp0_i_writemaster1_data_model_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:307:34  */
  assign dp0_i_n2612 = dp0_i_writemaster1_thread_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:312:31  */
  assign dp0_i_n2613 = dp0_i_readmaster2_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:313:31  */
  assign dp0_i_n2614 = dp0_i_readmaster2_fork_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:314:29  */
  assign dp0_i_n2615 = dp0_i_readmaster2_cs_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:315:31  */
  assign dp0_i_n2616 = dp0_i_readmaster2_read_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:316:34  */
  assign dp0_i_n2617 = dp0_i_readmaster2_read_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:317:38  */
  assign dp0_i_n2618 = dp0_i_readmaster2_read_vector_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:318:39  */
  assign dp0_i_n2619 = dp0_i_readmaster2_read_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:323:35  */
  assign dp0_i_n2620 = dp0_i_readmaster2_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:324:33  */
  assign dp0_i_n2621 = dp0_i_readmaster2_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:328:32  */
  assign dp0_i_n2622 = dp0_i_writemaster2_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:329:32  */
  assign dp0_i_n2623 = dp0_i_writemaster2_fork_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:330:30  */
  assign dp0_i_n2624 = dp0_i_writemaster2_cs_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:331:33  */
  assign dp0_i_n2625 = dp0_i_writemaster2_write_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:332:30  */
  assign dp0_i_n2626 = dp0_i_writemaster2_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:333:40  */
  assign dp0_i_n2627 = dp0_i_writemaster2_write_vector_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:334:41  */
  assign dp0_i_n2628 = dp0_i_writemaster2_write_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:335:37  */
  assign dp0_i_n2629 = dp0_i_writemaster2_writedata_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:337:36  */
  assign dp0_i_n2630 = dp0_i_writemaster2_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:338:34  */
  assign dp0_i_n2631 = dp0_i_writemaster2_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:339:34  */
  assign dp0_i_n2632 = dp0_i_writemaster2_thread_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:344:31  */
  assign dp0_i_n2633 = dp0_i_readmaster3_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:345:29  */
  assign dp0_i_n2634 = dp0_i_readmaster3_cs_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:346:31  */
  assign dp0_i_n2635 = dp0_i_readmaster3_read_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:347:34  */
  assign dp0_i_n2636 = dp0_i_readmaster3_read_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:348:38  */
  assign dp0_i_n2637 = dp0_i_readmaster3_read_vector_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:349:39  */
  assign dp0_i_n2638 = dp0_i_readmaster3_read_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:350:37  */
  assign dp0_i_n2639 = dp0_i_readmaster3_read_start_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:351:35  */
  assign dp0_i_n2640 = dp0_i_readmaster3_read_end_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:356:35  */
  assign dp0_i_n2641 = dp0_i_readmaster3_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:357:33  */
  assign dp0_i_n2642 = dp0_i_readmaster3_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:358:38  */
  assign dp0_i_n2643 = dp0_i_readmaster3_filler_data_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:362:32  */
  assign dp0_i_n2644 = dp0_i_writemaster3_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:363:30  */
  assign dp0_i_n2645 = dp0_i_writemaster3_cs_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:364:33  */
  assign dp0_i_n2646 = dp0_i_writemaster3_write_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:365:30  */
  assign dp0_i_n2647 = dp0_i_writemaster3_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:366:40  */
  assign dp0_i_n2648 = dp0_i_writemaster3_write_vector_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:367:41  */
  assign dp0_i_n2649 = dp0_i_writemaster3_write_scatter_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:368:37  */
  assign dp0_i_n2650 = dp0_i_writemaster3_write_end_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:369:37  */
  assign dp0_i_n2651 = dp0_i_writemaster3_writedata_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:371:36  */
  assign dp0_i_n2652 = dp0_i_writemaster3_burstlen_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:372:37  */
  assign dp0_i_n2653 = dp0_i_writemaster3_burstlen2_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:373:37  */
  assign dp0_i_n2654 = dp0_i_writemaster3_burstlen3_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:374:34  */
  assign dp0_i_n2655 = dp0_i_writemaster3_bus_id_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:375:34  */
  assign dp0_i_n2656 = dp0_i_writemaster3_thread_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:380:30  */
  assign dp0_i_n2657 = dp0_i_task_start_addr_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:381:19  */
  assign dp0_i_n2658 = dp0_i_task_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:383:22  */
  assign dp0_i_n2660 = dp0_i_task_vm_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:384:25  */
  assign dp0_i_n2661 = dp0_i_task_pcore_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:385:28  */
  assign dp0_i_n2662 = dp0_i_task_lockstep_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:386:28  */
  assign dp0_i_n2663 = dp0_i_task_tid_mask_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:387:34  */
  assign dp0_i_n2664 = dp0_i_task_iregister_auto_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:388:30  */
  assign dp0_i_n2665 = dp0_i_task_data_model_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:396:33  */
  assign dp0_i_n2666 = dp0_i_indication_avail_out; // (signal)
  /* ../../HW/src/dp/dp_core.vhd:238:1  */
  dp_0_611cf22eded7b64824a5f5c8e04751a6c8c2392b dp0_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .bus_waddr_in(bus_waddr_in),
    .bus_raddr_in(bus_raddr_in),
    .bus_write_in(bus_write_in),
    .bus_read_in(bus_read_in),
    .bus_writedata_in(bus_writedata_in),
    .readmaster1_readdatavalid_in(readmaster1_readdatavalid_in),
    .readmaster1_readdatavalid_vm_in(readmaster1_readdatavalid_vm_in),
    .readmaster1_readdata_in(readmaster1_readdata_in),
    .readmaster1_wait_request_in(readmaster1_wait_request_in),
    .writemaster1_wait_request_in(writemaster1_wait_request_in),
    .writemaster1_counter_in(writemaster1_counter_in),
    .readmaster2_readdatavalid_in(readmaster2_readdatavalid_in),
    .readmaster2_readdatavalid_vm_in(readmaster2_readdatavalid_vm_in),
    .readmaster2_readdata_in(readmaster2_readdata_in),
    .readmaster2_wait_request_in(readmaster2_wait_request_in),
    .writemaster2_wait_request_in(writemaster2_wait_request_in),
    .writemaster2_counter_in(writemaster2_counter_in),
    .readmaster3_readdatavalid_in(readmaster3_readdatavalid_in),
    .readmaster3_readdatavalid_vm_in(readmaster3_readdatavalid_vm_in),
    .readmaster3_readdata_in(readmaster3_readdata_in),
    .readmaster3_wait_request_in(readmaster3_wait_request_in),
    .writemaster3_wait_request_in(writemaster3_wait_request_in),
    .writemaster3_counter_in(writemaster3_counter_in),
    .task_busy_in(task_busy),
    .task_ready_in(task_ready),
    .bar_in(bar_in),
    .ddr_tx_busy_in(ddr_tx_busy_in),
    .bus_readdata_out(dp0_i_bus_readdata_out),
    .bus_readdatavalid_out(dp0_i_bus_readdatavalid_out),
    .bus_writewait_out(dp0_i_bus_writewait_out),
    .bus_readwait_out(dp0_i_bus_readwait_out),
    .readmaster1_addr_out(dp0_i_readmaster1_addr_out),
    .readmaster1_fork_out(dp0_i_readmaster1_fork_out),
    .readmaster1_addr_mode_out(dp0_i_readmaster1_addr_mode_out),
    .readmaster1_cs_out(dp0_i_readmaster1_cs_out),
    .readmaster1_read_out(dp0_i_readmaster1_read_out),
    .readmaster1_read_vm_out(dp0_i_readmaster1_read_vm_out),
    .readmaster1_read_data_flow_out(dp0_i_readmaster1_read_data_flow_out),
    .readmaster1_read_stream_out(dp0_i_readmaster1_read_stream_out),
    .readmaster1_read_stream_id_out(dp0_i_readmaster1_read_stream_id_out),
    .readmaster1_read_vector_out(dp0_i_readmaster1_read_vector_out),
    .readmaster1_read_scatter_out(dp0_i_readmaster1_read_scatter_out),
    .readmaster1_burstlen_out(dp0_i_readmaster1_burstlen_out),
    .readmaster1_bus_id_out(dp0_i_readmaster1_bus_id_out),
    .readmaster1_data_type_out(dp0_i_readmaster1_data_type_out),
    .readmaster1_data_model_out(dp0_i_readmaster1_data_model_out),
    .writemaster1_addr_out(dp0_i_writemaster1_addr_out),
    .writemaster1_fork_out(dp0_i_writemaster1_fork_out),
    .writemaster1_addr_mode_out(dp0_i_writemaster1_addr_mode_out),
    .writemaster1_vm_out(dp0_i_writemaster1_vm_out),
    .writemaster1_mcast_out(dp0_i_writemaster1_mcast_out),
    .writemaster1_cs_out(dp0_i_writemaster1_cs_out),
    .writemaster1_write_out(dp0_i_writemaster1_write_out),
    .writemaster1_write_data_flow_out(dp0_i_writemaster1_write_data_flow_out),
    .writemaster1_write_vector_out(dp0_i_writemaster1_write_vector_out),
    .writemaster1_write_stream_out(dp0_i_writemaster1_write_stream_out),
    .writemaster1_write_stream_id_out(dp0_i_writemaster1_write_stream_id_out),
    .writemaster1_write_scatter_out(dp0_i_writemaster1_write_scatter_out),
    .writemaster1_writedata_out(dp0_i_writemaster1_writedata_out),
    .writemaster1_burstlen_out(dp0_i_writemaster1_burstlen_out),
    .writemaster1_bus_id_out(dp0_i_writemaster1_bus_id_out),
    .writemaster1_data_type_out(dp0_i_writemaster1_data_type_out),
    .writemaster1_data_model_out(dp0_i_writemaster1_data_model_out),
    .writemaster1_thread_out(dp0_i_writemaster1_thread_out),
    .readmaster2_addr_out(dp0_i_readmaster2_addr_out),
    .readmaster2_fork_out(dp0_i_readmaster2_fork_out),
    .readmaster2_cs_out(dp0_i_readmaster2_cs_out),
    .readmaster2_read_out(dp0_i_readmaster2_read_out),
    .readmaster2_read_vm_out(dp0_i_readmaster2_read_vm_out),
    .readmaster2_read_vector_out(dp0_i_readmaster2_read_vector_out),
    .readmaster2_read_scatter_out(dp0_i_readmaster2_read_scatter_out),
    .readmaster2_burstlen_out(dp0_i_readmaster2_burstlen_out),
    .readmaster2_bus_id_out(dp0_i_readmaster2_bus_id_out),
    .writemaster2_addr_out(dp0_i_writemaster2_addr_out),
    .writemaster2_vm_out(dp0_i_writemaster2_vm_out),
    .writemaster2_fork_out(dp0_i_writemaster2_fork_out),
    .writemaster2_cs_out(dp0_i_writemaster2_cs_out),
    .writemaster2_write_out(dp0_i_writemaster2_write_out),
    .writemaster2_write_vector_out(dp0_i_writemaster2_write_vector_out),
    .writemaster2_write_scatter_out(dp0_i_writemaster2_write_scatter_out),
    .writemaster2_writedata_out(dp0_i_writemaster2_writedata_out),
    .writemaster2_burstlen_out(dp0_i_writemaster2_burstlen_out),
    .writemaster2_bus_id_out(dp0_i_writemaster2_bus_id_out),
    .writemaster2_thread_out(dp0_i_writemaster2_thread_out),
    .readmaster3_addr_out(dp0_i_readmaster3_addr_out),
    .readmaster3_cs_out(dp0_i_readmaster3_cs_out),
    .readmaster3_read_out(dp0_i_readmaster3_read_out),
    .readmaster3_read_vm_out(dp0_i_readmaster3_read_vm_out),
    .readmaster3_read_vector_out(dp0_i_readmaster3_read_vector_out),
    .readmaster3_read_scatter_out(dp0_i_readmaster3_read_scatter_out),
    .readmaster3_read_start_out(dp0_i_readmaster3_read_start_out),
    .readmaster3_read_end_out(dp0_i_readmaster3_read_end_out),
    .readmaster3_burstlen_out(dp0_i_readmaster3_burstlen_out),
    .readmaster3_bus_id_out(dp0_i_readmaster3_bus_id_out),
    .readmaster3_filler_data_out(dp0_i_readmaster3_filler_data_out),
    .writemaster3_addr_out(dp0_i_writemaster3_addr_out),
    .writemaster3_cs_out(dp0_i_writemaster3_cs_out),
    .writemaster3_write_out(dp0_i_writemaster3_write_out),
    .writemaster3_vm_out(dp0_i_writemaster3_vm_out),
    .writemaster3_write_vector_out(dp0_i_writemaster3_write_vector_out),
    .writemaster3_write_scatter_out(dp0_i_writemaster3_write_scatter_out),
    .writemaster3_write_end_out(dp0_i_writemaster3_write_end_out),
    .writemaster3_writedata_out(dp0_i_writemaster3_writedata_out),
    .writemaster3_burstlen_out(dp0_i_writemaster3_burstlen_out),
    .writemaster3_burstlen2_out(dp0_i_writemaster3_burstlen2_out),
    .writemaster3_burstlen3_out(dp0_i_writemaster3_burstlen3_out),
    .writemaster3_bus_id_out(dp0_i_writemaster3_bus_id_out),
    .writemaster3_thread_out(dp0_i_writemaster3_thread_out),
    .task_start_addr_out(dp0_i_task_start_addr_out),
    .task_out(dp0_i_task_out),
    .task_pending_out(),
    .task_vm_out(dp0_i_task_vm_out),
    .task_pcore_out(dp0_i_task_pcore_out),
    .task_lockstep_out(dp0_i_task_lockstep_out),
    .task_tid_mask_out(dp0_i_task_tid_mask_out),
    .task_iregister_auto_out(dp0_i_task_iregister_auto_out),
    .task_data_model_out(dp0_i_task_data_model_out),
    .indication_avail_out(dp0_i_indication_avail_out));
  /* ../../HW/src/dp/dp_core.vhd:408:40  */
  assign n2850_o = task_busy_in[0];
  /* ../../HW/src/dp/dp_core.vhd:408:49  */
  assign n2851_o = n2850_o | task_0_busy_r;
  /* ../../HW/src/dp/dp_core.vhd:408:21  */
  assign n2852_o = n2851_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_core.vhd:412:40  */
  assign n2855_o = task_busy_in[1];
  /* ../../HW/src/dp/dp_core.vhd:412:49  */
  assign n2856_o = n2855_o | task_1_busy_r;
  /* ../../HW/src/dp/dp_core.vhd:412:21  */
  assign n2857_o = n2856_o ? 1'b1 : 1'b0;
  /* ../../HW/src/dp/dp_core.vhd:416:41  */
  assign n2860_o = ~task_ready_in;
  /* ../../HW/src/dp/dp_core.vhd:416:47  */
  assign n2861_o = n2860_o | task_busy_r;
  /* ../../HW/src/dp/dp_core.vhd:416:21  */
  assign n2862_o = n2861_o ? 1'b0 : 1'b1;
  /* ../../HW/src/dp/dp_core.vhd:429:13  */
  assign n2866_o = ~reset_in;
  /* ../../HW/src/dp/dp_core.vhd:472:38  */
  assign n2868_o = task_rrrrrrrr | task_rrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:473:37  */
  assign n2869_o = n2868_o | task_rrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:474:36  */
  assign n2870_o = n2869_o | task_rrrrr;
  /* ../../HW/src/dp/dp_core.vhd:475:35  */
  assign n2871_o = n2870_o | task_rrrr;
  /* ../../HW/src/dp/dp_core.vhd:476:34  */
  assign n2872_o = n2871_o | task_rrr;
  /* ../../HW/src/dp/dp_core.vhd:477:33  */
  assign n2873_o = n2872_o | task_rr;
  /* ../../HW/src/dp/dp_core.vhd:478:32  */
  assign n2874_o = n2873_o | task_r;
  /* ../../HW/src/dp/dp_core.vhd:479:31  */
  assign n2875_o = n2874_o | \task ;
  /* ../../HW/src/dp/dp_core.vhd:482:46  */
  assign n2876_o = ~task_vm_rrrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:482:41  */
  assign n2877_o = task_rrrrrrrr & n2876_o;
  /* ../../HW/src/dp/dp_core.vhd:483:37  */
  assign n2878_o = ~task_vm_rrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:483:32  */
  assign n2879_o = task_rrrrrrr & n2878_o;
  /* ../../HW/src/dp/dp_core.vhd:482:69  */
  assign n2880_o = n2877_o | n2879_o;
  /* ../../HW/src/dp/dp_core.vhd:484:36  */
  assign n2881_o = ~task_vm_rrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:484:31  */
  assign n2882_o = task_rrrrrr & n2881_o;
  /* ../../HW/src/dp/dp_core.vhd:483:59  */
  assign n2883_o = n2880_o | n2882_o;
  /* ../../HW/src/dp/dp_core.vhd:485:35  */
  assign n2884_o = ~task_vm_rrrrr;
  /* ../../HW/src/dp/dp_core.vhd:485:30  */
  assign n2885_o = task_rrrrr & n2884_o;
  /* ../../HW/src/dp/dp_core.vhd:484:57  */
  assign n2886_o = n2883_o | n2885_o;
  /* ../../HW/src/dp/dp_core.vhd:486:42  */
  assign n2887_o = ~task_vm_rrrr;
  /* ../../HW/src/dp/dp_core.vhd:486:37  */
  assign n2888_o = task_rrrr & n2887_o;
  /* ../../HW/src/dp/dp_core.vhd:485:55  */
  assign n2889_o = n2886_o | n2888_o;
  /* ../../HW/src/dp/dp_core.vhd:487:33  */
  assign n2890_o = ~task_vm_rrr;
  /* ../../HW/src/dp/dp_core.vhd:487:28  */
  assign n2891_o = task_rrr & n2890_o;
  /* ../../HW/src/dp/dp_core.vhd:486:61  */
  assign n2892_o = n2889_o | n2891_o;
  /* ../../HW/src/dp/dp_core.vhd:488:40  */
  assign n2893_o = ~task_vm_rr;
  /* ../../HW/src/dp/dp_core.vhd:488:35  */
  assign n2894_o = task_rr & n2893_o;
  /* ../../HW/src/dp/dp_core.vhd:487:51  */
  assign n2895_o = n2892_o | n2894_o;
  /* ../../HW/src/dp/dp_core.vhd:489:39  */
  assign n2896_o = ~task_vm_r;
  /* ../../HW/src/dp/dp_core.vhd:489:34  */
  assign n2897_o = task_r & n2896_o;
  /* ../../HW/src/dp/dp_core.vhd:488:57  */
  assign n2898_o = n2895_o | n2897_o;
  /* ../../HW/src/dp/dp_core.vhd:490:37  */
  assign n2899_o = ~task_vm;
  /* ../../HW/src/dp/dp_core.vhd:490:32  */
  assign n2900_o = \task  & n2899_o;
  /* ../../HW/src/dp/dp_core.vhd:489:55  */
  assign n2901_o = n2898_o | n2900_o;
  /* ../../HW/src/dp/dp_core.vhd:493:41  */
  assign n2902_o = task_rrrrrrrr & task_vm_rrrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:494:32  */
  assign n2903_o = task_rrrrrrr & task_vm_rrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:493:65  */
  assign n2904_o = n2902_o | n2903_o;
  /* ../../HW/src/dp/dp_core.vhd:495:31  */
  assign n2905_o = task_rrrrrr & task_vm_rrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:494:55  */
  assign n2906_o = n2904_o | n2905_o;
  /* ../../HW/src/dp/dp_core.vhd:496:30  */
  assign n2907_o = task_rrrrr & task_vm_rrrrr;
  /* ../../HW/src/dp/dp_core.vhd:495:53  */
  assign n2908_o = n2906_o | n2907_o;
  /* ../../HW/src/dp/dp_core.vhd:497:37  */
  assign n2909_o = task_rrrr & task_vm_rrrr;
  /* ../../HW/src/dp/dp_core.vhd:496:51  */
  assign n2910_o = n2908_o | n2909_o;
  /* ../../HW/src/dp/dp_core.vhd:498:36  */
  assign n2911_o = task_rrr & task_vm_rrr;
  /* ../../HW/src/dp/dp_core.vhd:497:57  */
  assign n2912_o = n2910_o | n2911_o;
  /* ../../HW/src/dp/dp_core.vhd:499:35  */
  assign n2913_o = task_rr & task_vm_rr;
  /* ../../HW/src/dp/dp_core.vhd:498:55  */
  assign n2914_o = n2912_o | n2913_o;
  /* ../../HW/src/dp/dp_core.vhd:500:34  */
  assign n2915_o = task_r & task_vm_r;
  /* ../../HW/src/dp/dp_core.vhd:499:53  */
  assign n2916_o = n2914_o | n2915_o;
  /* ../../HW/src/dp/dp_core.vhd:501:32  */
  assign n2917_o = \task  & task_vm;
  /* ../../HW/src/dp/dp_core.vhd:500:51  */
  assign n2918_o = n2916_o | n2917_o;
  assign n2995_o = {n2857_o, n2852_o};
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n2996_q <= 5'b11111;
    else
      n2996_q <= task_pcore;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n2997_q <= 1'b0;
    else
      n2997_q <= task_lockstep;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n2998_q <= 4'b0000;
    else
      n2998_q <= task_tid_mask;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n2999_q <= 28'b0000000000000000000000000000;
    else
      n2999_q <= task_iregister_auto;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3000_q <= 2'b00;
    else
      n3000_q <= task_data_model;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3001_q <= 11'b00000000000;
    else
      n3001_q <= task_start_addr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3002_q <= 1'b0;
    else
      n3002_q <= \task ;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3003_q <= 1'b0;
    else
      n3003_q <= task_r;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3004_q <= 1'b0;
    else
      n3004_q <= task_rr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3005_q <= 1'b0;
    else
      n3005_q <= task_rrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3006_q <= 1'b0;
    else
      n3006_q <= task_rrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3007_q <= 1'b0;
    else
      n3007_q <= task_rrrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3008_q <= 1'b0;
    else
      n3008_q <= task_rrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3009_q <= 1'b0;
    else
      n3009_q <= task_rrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3010_q <= 1'b0;
    else
      n3010_q <= task_vm;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3011_q <= 1'b0;
    else
      n3011_q <= task_vm_r;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3012_q <= 1'b0;
    else
      n3012_q <= task_vm_rr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3013_q <= 1'b0;
    else
      n3013_q <= task_vm_rrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3014_q <= 1'b0;
    else
      n3014_q <= task_vm_rrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3015_q <= 1'b0;
    else
      n3015_q <= task_vm_rrrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3016_q <= 1'b0;
    else
      n3016_q <= task_vm_rrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3017_q <= 1'b0;
    else
      n3017_q <= task_vm_rrrrrrr;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3018_q <= 1'b0;
    else
      n3018_q <= n2875_o;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3019_q <= 1'b0;
    else
      n3019_q <= n2918_o;
  /* ../../HW/src/dp/dp_core.vhd:456:5  */
  always @(posedge clock_in or posedge n2866_o)
    if (n2866_o)
      n3020_q <= 1'b0;
    else
      n3020_q <= n2901_o;
endmodule

module ddr_tx
  (input  clock_in,
   input  reset_in,
   input  [31:0] write_addr_in,
   input  write_cs_in,
   input  write_in,
   input  [2:0] write_vector_in,
   input  [3:0] write_end_in,
   input  [63:0] write_data_in,
   input  [4:0] write_burstlen_in,
   input  [8:0] write_burstlen2_in,
   input  [4:0] write_burstlen3_in,
   input  ddr_awready_in,
   input  ddr_wready_in,
   input  ddr_bresp_in,
   output write_wait_request_out,
   output [31:0] ddr_awaddr_out,
   output [2:0] ddr_awlen_out,
   output ddr_awvalid_out,
   output [31:0] ddr_waddr_out,
   output ddr_wvalid_out,
   output [63:0] ddr_wdata_out,
   output ddr_wlast_out,
   output [7:0] ddr_wbe_out,
   output [1:0] ddr_awburst_out,
   output [3:0] ddr_awcache_out,
   output ddr_awid_out,
   output ddr_awlock_out,
   output [2:0] ddr_awprot_out,
   output [3:0] ddr_awqos_out,
   output [2:0] ddr_awsize_out,
   output ddr_bready_out,
   output ddr_tx_busy_out);
  wire write2;
  wire ddr_write;
  wire [15:0] byteenable;
  wire [40:0] write_data_write_r;
  wire [40:0] write_data_write;
  wire write_data_write_ena;
  wire write_data_write_ena_r;
  wire [127:0] write_data;
  wire [127:0] write_data_r;
  wire [63:0] write_data_2_r;
  wire [15:0] byteenable_r;
  wire [31:0] wr_ddr_addr;
  wire [31:0] write_next_addr_r;
  wire w_x1;
  wire w_x2;
  wire w_x4;
  wire w_x8;
  wire w_mask1;
  wire w_mask2;
  wire w_mask3;
  wire w_mask4;
  wire w_mask5;
  wire w_mask6;
  wire w_mask7;
  wire w_mask8;
  wire write_complete;
  wire write_over_complete;
  wire write_flush_r;
  wire [9:0] write_request_r;
  wire [9:0] write_complete_r;
  wire ready;
  wire hold;
  wire awvalid;
  wire [2:0] awlen_r;
  wire [31:0] awaddr_r;
  wire n1572_o;
  wire n1573_o;
  wire n1574_o;
  wire n1575_o;
  wire [31:0] n1576_o;
  wire n1578_o;
  wire [31:0] n1579_o;
  wire [31:0] n1580_o;
  wire [7:0] n1581_o;
  localparam [1:0] n1582_o = 2'b01;
  localparam [3:0] n1583_o = 4'b0011;
  localparam n1584_o = 1'b0;
  localparam n1585_o = 1'b0;
  localparam [2:0] n1586_o = 3'b000;
  localparam [3:0] n1587_o = 4'b0000;
  localparam n1588_o = 1'b1;
  localparam [2:0] n1589_o = 3'b011;
  wire n1591_o;
  wire n1592_o;
  wire n1593_o;
  wire n1594_o;
  wire [2:0] n1597_o;
  wire [3:0] n1599_o;
  wire [3:0] n1601_o;
  wire [3:0] n1602_o;
  wire [3:0] n1604_o;
  wire n1606_o;
  wire n1607_o;
  wire [2:0] n1610_o;
  wire [3:0] n1612_o;
  wire [3:0] n1614_o;
  wire [3:0] n1615_o;
  wire [3:0] n1617_o;
  wire n1619_o;
  wire n1620_o;
  wire n1624_o;
  wire n1625_o;
  wire n1626_o;
  wire n1627_o;
  wire n1628_o;
  wire n1629_o;
  wire n1630_o;
  wire n1632_o;
  wire n1634_o;
  wire n1635_o;
  wire n1636_o;
  wire n1637_o;
  wire n1638_o;
  wire n1641_o;
  wire n1642_o;
  wire n1645_o;
  wire n1647_o;
  wire n1648_o;
  wire n1649_o;
  wire n1650_o;
  wire n1654_o;
  wire n1657_o;
  wire n1658_o;
  wire [31:0] n1659_o;
  wire [9:0] n1662_o;
  wire [2:0] n1664_o;
  wire [2:0] n1665_o;
  wire [2:0] n1668_o;
  wire n1681_o;
  wire [7:0] n1682_o;
  wire [31:0] n1683_o;
  wire n1685_o;
  wire n1688_o;
  wire [7:0] n1689_o;
  wire [40:0] n1691_o;
  wire [40:0] n1692_o;
  wire [40:0] n1693_o;
  wire [28:0] n1698_o;
  wire [31:0] n1700_o;
  wire n1705_o;
  wire n1707_o;
  wire n1709_o;
  wire n1711_o;
  wire n1712_o;
  wire n1715_o;
  wire n1717_o;
  wire [31:0] n1720_o;
  wire [9:0] n1723_o;
  wire n1741_o;
  wire n1743_o;
  wire n1745_o;
  wire n1748_o;
  wire n1751_o;
  wire n1754_o;
  wire n1756_o;
  wire n1758_o;
  wire n1760_o;
  wire n1762_o;
  wire n1764_o;
  wire n1766_o;
  wire n1771_o;
  wire n1772_o;
  wire n1776_o;
  wire n1777_o;
  wire n1781_o;
  wire n1782_o;
  wire n1786_o;
  wire n1787_o;
  wire n1791_o;
  wire n1792_o;
  wire n1796_o;
  wire n1797_o;
  wire n1801_o;
  wire n1802_o;
  wire n1806_o;
  wire n1807_o;
  wire [2:0] n1811_o;
  wire n1812_o;
  wire n1813_o;
  wire n1814_o;
  wire n1815_o;
  wire n1816_o;
  wire n1817_o;
  wire n1818_o;
  wire n1819_o;
  wire n1820_o;
  wire n1821_o;
  wire n1822_o;
  wire n1823_o;
  wire n1824_o;
  wire n1825_o;
  wire n1826_o;
  wire n1827_o;
  wire n1828_o;
  wire n1829_o;
  wire n1830_o;
  wire n1831_o;
  wire n1832_o;
  wire n1833_o;
  wire n1834_o;
  wire n1835_o;
  wire n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire n1843_o;
  wire n1845_o;
  wire n1846_o;
  wire n1847_o;
  wire n1848_o;
  wire n1849_o;
  wire n1850_o;
  wire n1851_o;
  wire n1852_o;
  wire n1853_o;
  wire n1854_o;
  wire n1855_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1859_o;
  wire n1860_o;
  wire n1861_o;
  wire n1862_o;
  wire n1863_o;
  wire n1864_o;
  wire n1865_o;
  wire n1866_o;
  wire n1867_o;
  wire n1868_o;
  wire n1869_o;
  wire n1870_o;
  wire n1871_o;
  wire n1872_o;
  wire n1873_o;
  wire n1874_o;
  wire n1875_o;
  wire n1876_o;
  wire n1877_o;
  wire n1879_o;
  wire n1880_o;
  wire n1881_o;
  wire n1882_o;
  wire n1883_o;
  wire n1884_o;
  wire n1885_o;
  wire n1886_o;
  wire n1887_o;
  wire n1888_o;
  wire n1889_o;
  wire n1890_o;
  wire n1891_o;
  wire n1892_o;
  wire n1893_o;
  wire n1894_o;
  wire n1895_o;
  wire n1896_o;
  wire n1897_o;
  wire n1898_o;
  wire n1899_o;
  wire n1900_o;
  wire n1901_o;
  wire n1902_o;
  wire n1903_o;
  wire n1904_o;
  wire n1905_o;
  wire n1906_o;
  wire n1907_o;
  wire n1908_o;
  wire n1909_o;
  wire n1910_o;
  wire n1911_o;
  wire n1913_o;
  wire n1914_o;
  wire n1915_o;
  wire n1916_o;
  wire n1917_o;
  wire n1918_o;
  wire n1919_o;
  wire n1920_o;
  wire n1921_o;
  wire n1922_o;
  wire n1923_o;
  wire n1924_o;
  wire n1925_o;
  wire n1926_o;
  wire n1927_o;
  wire n1928_o;
  wire n1929_o;
  wire n1930_o;
  wire n1931_o;
  wire n1932_o;
  wire n1933_o;
  wire n1934_o;
  wire n1935_o;
  wire n1936_o;
  wire n1937_o;
  wire n1938_o;
  wire n1939_o;
  wire n1940_o;
  wire n1941_o;
  wire n1942_o;
  wire n1943_o;
  wire n1944_o;
  wire n1945_o;
  wire n1947_o;
  wire n1948_o;
  wire n1949_o;
  wire n1950_o;
  wire n1951_o;
  wire n1952_o;
  wire n1953_o;
  wire n1954_o;
  wire n1955_o;
  wire n1956_o;
  wire n1957_o;
  wire n1958_o;
  wire n1959_o;
  wire n1960_o;
  wire n1961_o;
  wire n1962_o;
  wire n1963_o;
  wire n1964_o;
  wire n1965_o;
  wire n1966_o;
  wire n1967_o;
  wire n1968_o;
  wire n1969_o;
  wire n1970_o;
  wire n1971_o;
  wire n1972_o;
  wire n1973_o;
  wire n1974_o;
  wire n1975_o;
  wire n1976_o;
  wire n1977_o;
  wire n1978_o;
  wire n1979_o;
  wire n1981_o;
  wire n1982_o;
  wire n1983_o;
  wire n1984_o;
  wire n1985_o;
  wire n1986_o;
  wire n1987_o;
  wire n1988_o;
  wire n1989_o;
  wire n1990_o;
  wire n1991_o;
  wire n1992_o;
  wire n1993_o;
  wire n1994_o;
  wire n1995_o;
  wire n1996_o;
  wire n1997_o;
  wire n1998_o;
  wire n1999_o;
  wire n2000_o;
  wire n2001_o;
  wire n2002_o;
  wire n2003_o;
  wire n2004_o;
  wire n2005_o;
  wire n2006_o;
  wire n2007_o;
  wire n2008_o;
  wire n2009_o;
  wire n2010_o;
  wire n2011_o;
  wire n2012_o;
  wire n2013_o;
  wire n2015_o;
  wire n2016_o;
  wire n2017_o;
  wire n2018_o;
  wire n2019_o;
  wire n2020_o;
  wire n2021_o;
  wire n2022_o;
  wire n2023_o;
  wire n2024_o;
  wire n2025_o;
  wire n2026_o;
  wire n2027_o;
  wire n2028_o;
  wire n2029_o;
  wire n2030_o;
  wire n2031_o;
  wire n2032_o;
  wire n2033_o;
  wire n2034_o;
  wire n2035_o;
  wire n2036_o;
  wire n2037_o;
  wire n2038_o;
  wire n2039_o;
  wire n2040_o;
  wire n2041_o;
  wire n2042_o;
  wire n2043_o;
  wire n2044_o;
  wire n2045_o;
  wire n2046_o;
  wire n2047_o;
  wire n2049_o;
  wire n2050_o;
  wire n2051_o;
  wire n2052_o;
  wire n2053_o;
  wire n2054_o;
  wire n2055_o;
  wire n2056_o;
  wire n2057_o;
  wire n2058_o;
  wire n2059_o;
  wire n2060_o;
  wire n2061_o;
  wire n2062_o;
  wire n2063_o;
  wire n2064_o;
  wire n2065_o;
  wire n2066_o;
  wire n2067_o;
  wire n2068_o;
  wire n2069_o;
  wire n2070_o;
  wire n2071_o;
  wire n2072_o;
  wire n2073_o;
  wire n2074_o;
  wire n2075_o;
  wire n2076_o;
  wire n2077_o;
  wire n2078_o;
  wire n2079_o;
  wire n2080_o;
  wire n2081_o;
  wire [6:0] n2082_o;
  reg n2083_o;
  reg n2084_o;
  reg n2085_o;
  reg n2086_o;
  reg n2087_o;
  reg n2088_o;
  reg n2089_o;
  reg n2090_o;
  reg n2091_o;
  reg n2092_o;
  reg n2093_o;
  reg n2094_o;
  reg n2095_o;
  reg n2096_o;
  reg n2097_o;
  reg n2098_o;
  wire [15:0] n2099_o;
  wire [15:0] n2100_o;
  wire [2:0] n2104_o;
  wire n2106_o;
  wire [31:0] n2107_o;
  wire n2109_o;
  wire [15:0] n2110_o;
  wire n2112_o;
  wire [7:0] n2113_o;
  wire [7:0] n2114_o;
  wire [7:0] n2115_o;
  wire [55:0] n2116_o;
  wire [55:0] n2117_o;
  wire [55:0] n2118_o;
  wire [63:0] n2119_o;
  wire [15:0] n2120_o;
  wire [15:0] n2121_o;
  wire [47:0] n2122_o;
  wire [47:0] n2123_o;
  wire [47:0] n2124_o;
  wire [63:0] n2125_o;
  wire [31:0] n2126_o;
  wire [31:0] n2127_o;
  wire [31:0] n2128_o;
  wire [31:0] n2129_o;
  wire [31:0] n2130_o;
  wire n2132_o;
  wire n2134_o;
  wire [31:0] n2135_o;
  wire n2137_o;
  wire [15:0] n2138_o;
  wire n2140_o;
  wire [7:0] n2141_o;
  wire [7:0] n2142_o;
  wire [7:0] n2143_o;
  wire [55:0] n2144_o;
  wire [55:0] n2145_o;
  wire [55:0] n2146_o;
  wire [63:0] n2147_o;
  wire [15:0] n2148_o;
  wire [15:0] n2149_o;
  wire [47:0] n2150_o;
  wire [47:0] n2151_o;
  wire [47:0] n2152_o;
  wire [63:0] n2153_o;
  wire [31:0] n2154_o;
  wire [31:0] n2155_o;
  wire [31:0] n2156_o;
  wire [31:0] n2157_o;
  wire [31:0] n2158_o;
  wire n2160_o;
  wire n2162_o;
  wire [31:0] n2163_o;
  wire n2165_o;
  wire [15:0] n2166_o;
  wire n2168_o;
  wire [7:0] n2169_o;
  wire [7:0] n2170_o;
  wire [7:0] n2171_o;
  wire [55:0] n2172_o;
  wire [55:0] n2173_o;
  wire [55:0] n2174_o;
  wire [63:0] n2175_o;
  wire [15:0] n2176_o;
  wire [15:0] n2177_o;
  wire [47:0] n2178_o;
  wire [47:0] n2179_o;
  wire [47:0] n2180_o;
  wire [63:0] n2181_o;
  wire [31:0] n2182_o;
  wire [31:0] n2183_o;
  wire [31:0] n2184_o;
  wire [31:0] n2185_o;
  wire [31:0] n2186_o;
  wire n2188_o;
  wire n2190_o;
  wire [31:0] n2191_o;
  wire n2193_o;
  wire [15:0] n2194_o;
  wire n2196_o;
  wire [7:0] n2197_o;
  wire [7:0] n2198_o;
  wire [7:0] n2199_o;
  wire [55:0] n2200_o;
  wire [55:0] n2201_o;
  wire [55:0] n2202_o;
  wire [63:0] n2203_o;
  wire [15:0] n2204_o;
  wire [15:0] n2205_o;
  wire [47:0] n2206_o;
  wire [47:0] n2207_o;
  wire [47:0] n2208_o;
  wire [63:0] n2209_o;
  wire [31:0] n2210_o;
  wire [31:0] n2211_o;
  wire [31:0] n2212_o;
  wire [31:0] n2213_o;
  wire [31:0] n2214_o;
  wire n2216_o;
  wire n2218_o;
  wire [31:0] n2219_o;
  wire n2221_o;
  wire [15:0] n2222_o;
  wire n2224_o;
  wire [7:0] n2225_o;
  wire [7:0] n2226_o;
  wire [7:0] n2227_o;
  wire [55:0] n2228_o;
  wire [55:0] n2229_o;
  wire [55:0] n2230_o;
  wire [63:0] n2231_o;
  wire [15:0] n2232_o;
  wire [15:0] n2233_o;
  wire [47:0] n2234_o;
  wire [47:0] n2235_o;
  wire [47:0] n2236_o;
  wire [63:0] n2237_o;
  wire [31:0] n2238_o;
  wire [31:0] n2239_o;
  wire [31:0] n2240_o;
  wire [31:0] n2241_o;
  wire [31:0] n2242_o;
  wire n2244_o;
  wire n2246_o;
  wire [31:0] n2247_o;
  wire n2249_o;
  wire [15:0] n2250_o;
  wire n2252_o;
  wire [7:0] n2253_o;
  wire [7:0] n2254_o;
  wire [7:0] n2255_o;
  wire [55:0] n2256_o;
  wire [55:0] n2257_o;
  wire [55:0] n2258_o;
  wire [63:0] n2259_o;
  wire [15:0] n2260_o;
  wire [15:0] n2261_o;
  wire [47:0] n2262_o;
  wire [47:0] n2263_o;
  wire [47:0] n2264_o;
  wire [63:0] n2265_o;
  wire [31:0] n2266_o;
  wire [31:0] n2267_o;
  wire [31:0] n2268_o;
  wire [31:0] n2269_o;
  wire [31:0] n2270_o;
  wire n2272_o;
  wire n2274_o;
  wire [31:0] n2275_o;
  wire n2277_o;
  wire [15:0] n2278_o;
  wire n2280_o;
  wire [7:0] n2281_o;
  wire [7:0] n2282_o;
  wire [7:0] n2283_o;
  wire [55:0] n2284_o;
  wire [55:0] n2285_o;
  wire [55:0] n2286_o;
  wire [63:0] n2287_o;
  wire [15:0] n2288_o;
  wire [15:0] n2289_o;
  wire [47:0] n2290_o;
  wire [47:0] n2291_o;
  wire [47:0] n2292_o;
  wire [63:0] n2293_o;
  wire [31:0] n2294_o;
  wire [31:0] n2295_o;
  wire [31:0] n2296_o;
  wire [31:0] n2297_o;
  wire [31:0] n2298_o;
  wire n2300_o;
  wire n2302_o;
  wire [31:0] n2303_o;
  wire n2305_o;
  wire [15:0] n2306_o;
  wire n2308_o;
  wire [7:0] n2309_o;
  wire [7:0] n2310_o;
  wire [7:0] n2311_o;
  wire [55:0] n2312_o;
  wire [55:0] n2313_o;
  wire [55:0] n2314_o;
  wire [63:0] n2315_o;
  wire [15:0] n2316_o;
  wire [15:0] n2317_o;
  wire [47:0] n2318_o;
  wire [47:0] n2319_o;
  wire [47:0] n2320_o;
  wire [63:0] n2321_o;
  wire [31:0] n2322_o;
  wire [31:0] n2323_o;
  wire [31:0] n2324_o;
  wire [31:0] n2325_o;
  wire [31:0] n2326_o;
  wire [6:0] n2327_o;
  wire [7:0] n2328_o;
  wire [7:0] n2329_o;
  reg [7:0] n2330_o;
  wire [7:0] n2331_o;
  wire [7:0] n2332_o;
  wire [7:0] n2333_o;
  reg [7:0] n2334_o;
  wire [7:0] n2335_o;
  wire [7:0] n2336_o;
  wire [7:0] n2337_o;
  wire [7:0] n2338_o;
  reg [7:0] n2339_o;
  wire [7:0] n2340_o;
  wire [7:0] n2341_o;
  wire [7:0] n2342_o;
  wire [7:0] n2343_o;
  wire [7:0] n2344_o;
  reg [7:0] n2345_o;
  wire [7:0] n2346_o;
  wire [7:0] n2347_o;
  wire [7:0] n2348_o;
  wire [7:0] n2349_o;
  wire [7:0] n2350_o;
  wire [7:0] n2351_o;
  reg [7:0] n2352_o;
  wire [7:0] n2353_o;
  wire [7:0] n2354_o;
  wire [7:0] n2355_o;
  wire [7:0] n2356_o;
  wire [7:0] n2357_o;
  wire [7:0] n2358_o;
  wire [7:0] n2359_o;
  reg [7:0] n2360_o;
  wire [7:0] n2361_o;
  wire [7:0] n2362_o;
  wire [7:0] n2363_o;
  wire [7:0] n2364_o;
  wire [7:0] n2365_o;
  wire [7:0] n2366_o;
  wire [7:0] n2367_o;
  wire [7:0] n2368_o;
  reg [7:0] n2369_o;
  wire [7:0] n2370_o;
  wire [7:0] n2371_o;
  wire [7:0] n2372_o;
  wire [7:0] n2373_o;
  wire [7:0] n2374_o;
  wire [7:0] n2375_o;
  wire [7:0] n2376_o;
  wire [7:0] n2377_o;
  reg [7:0] n2378_o;
  wire [7:0] n2379_o;
  wire [7:0] n2380_o;
  wire [7:0] n2381_o;
  wire [7:0] n2382_o;
  wire [7:0] n2383_o;
  wire [7:0] n2384_o;
  wire [7:0] n2385_o;
  wire [7:0] n2386_o;
  reg [7:0] n2387_o;
  wire [7:0] n2388_o;
  wire [7:0] n2389_o;
  wire [7:0] n2390_o;
  wire [7:0] n2391_o;
  wire [7:0] n2392_o;
  wire [7:0] n2393_o;
  wire [7:0] n2394_o;
  reg [7:0] n2395_o;
  wire [7:0] n2396_o;
  wire [7:0] n2397_o;
  wire [7:0] n2398_o;
  wire [7:0] n2399_o;
  wire [7:0] n2400_o;
  wire [7:0] n2401_o;
  reg [7:0] n2402_o;
  wire [7:0] n2403_o;
  wire [7:0] n2404_o;
  wire [7:0] n2405_o;
  wire [7:0] n2406_o;
  wire [7:0] n2407_o;
  reg [7:0] n2408_o;
  wire [7:0] n2409_o;
  wire [7:0] n2410_o;
  wire [7:0] n2411_o;
  wire [7:0] n2412_o;
  reg [7:0] n2413_o;
  wire [7:0] n2414_o;
  wire [7:0] n2415_o;
  wire [7:0] n2416_o;
  reg [7:0] n2417_o;
  wire [7:0] n2418_o;
  wire [7:0] n2419_o;
  reg [7:0] n2420_o;
  wire [119:0] n2421_o;
  wire [119:0] n2422_o;
  wire [119:0] n2423_o;
  wire [7:0] n2424_o;
  wire n2428_o;
  wire [7:0] n2430_o;
  wire [63:0] n2432_o;
  wire [63:0] n2433_o;
  wire [127:0] n2434_o;
  wire [15:0] n2435_o;
  wire [63:0] n2437_o;
  wire [63:0] n2438_o;
  wire [63:0] n2439_o;
  wire [63:0] n2440_o;
  wire [63:0] n2441_o;
  wire [15:0] n2443_o;
  wire [15:0] n2444_o;
  wire [127:0] n2446_o;
  wire [40:0] n2459_o;
  reg [40:0] n2460_q;
  wire n2461_o;
  reg n2462_q;
  wire [127:0] n2466_o;
  reg [127:0] n2467_q;
  wire [63:0] n2468_o;
  reg [63:0] n2469_q;
  reg [15:0] n2470_q;
  wire [31:0] n2472_o;
  reg [31:0] n2473_q;
  wire n2474_o;
  reg n2475_q;
  wire [9:0] n2476_o;
  reg [9:0] n2477_q;
  wire [9:0] n2478_o;
  reg [9:0] n2479_q;
  reg [2:0] n2480_q;
  wire [31:0] n2481_o;
  reg [31:0] n2482_q;
  assign write_wait_request_out = n1642_o;
  assign ddr_awaddr_out = n1579_o;
  assign ddr_awlen_out = awlen_r;
  assign ddr_awvalid_out = awvalid;
  assign ddr_waddr_out = n1580_o;
  assign ddr_wvalid_out = ddr_write;
  assign ddr_wdata_out = write_data_2_r;
  assign ddr_wlast_out = awvalid;
  assign ddr_wbe_out = n1581_o;
  assign ddr_awburst_out = n1582_o;
  assign ddr_awcache_out = n1583_o;
  assign ddr_awid_out = n1584_o;
  assign ddr_awlock_out = n1585_o;
  assign ddr_awprot_out = n1586_o;
  assign ddr_awqos_out = n1587_o;
  assign ddr_awsize_out = n1589_o;
  assign ddr_bready_out = n1588_o;
  assign ddr_tx_busy_out = n1594_o;
  /* ../../HW/src/top/ddr_tx.vhd:99:8  */
  assign write2 = n1638_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:101:8  */
  assign ddr_write = n1575_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:102:8  */
  assign byteenable = n2100_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:103:8  */
  assign write_data_write_r = n2460_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:104:8  */
  assign write_data_write = n1693_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:105:8  */
  assign write_data_write_ena = n1630_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:106:8  */
  assign write_data_write_ena_r = n2462_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:110:8  */
  assign write_data = n2466_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:111:8  */
  assign write_data_r = n2467_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:112:8  */
  assign write_data_2_r = n2469_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:113:8  */
  assign byteenable_r = n2470_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:115:8  */
  assign wr_ddr_addr = n1700_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:116:8  */
  assign write_next_addr_r = n2473_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:118:8  */
  assign w_x1 = 1'b1; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:119:8  */
  assign w_x2 = n1762_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:120:8  */
  assign w_x4 = n1764_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:121:8  */
  assign w_x8 = n1766_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:123:8  */
  assign w_mask1 = n1772_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:124:8  */
  assign w_mask2 = n1777_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:125:8  */
  assign w_mask3 = n1782_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:126:8  */
  assign w_mask4 = n1787_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:127:8  */
  assign w_mask5 = n1792_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:128:8  */
  assign w_mask6 = n1797_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:129:8  */
  assign w_mask7 = n1802_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:130:8  */
  assign w_mask8 = n1807_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:132:8  */
  assign write_complete = n1607_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:133:8  */
  assign write_over_complete = n1620_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:134:8  */
  assign write_flush_r = n2475_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:136:8  */
  assign write_request_r = n2477_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:137:8  */
  assign write_complete_r = n2479_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:139:8  */
  assign ready = n1572_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:140:8  */
  assign hold = n1574_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:141:8  */
  assign awvalid = n1650_o; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:142:8  */
  assign awlen_r = n2480_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:143:8  */
  assign awaddr_r = n2482_q; // (signal)
  /* ../../HW/src/top/ddr_tx.vhd:152:25  */
  assign n1572_o = ddr_awready_in & ddr_wready_in;
  /* ../../HW/src/top/ddr_tx.vhd:154:37  */
  assign n1573_o = ~ready;
  /* ../../HW/src/top/ddr_tx.vhd:154:32  */
  assign n1574_o = write_data_write_ena_r & n1573_o;
  /* ../../HW/src/top/ddr_tx.vhd:156:37  */
  assign n1575_o = write_data_write_ena_r & ready;
  /* ../../HW/src/top/ddr_tx.vhd:162:38  */
  assign n1576_o = write_data_write_r[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:162:55  */
  assign n1578_o = awlen_r == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:162:43  */
  assign n1579_o = n1578_o ? n1576_o : awaddr_r;
  /* ../../HW/src/top/ddr_tx.vhd:170:37  */
  assign n1580_o = write_data_write_r[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:174:35  */
  assign n1581_o = write_data_write_r[39:32];
  /* ../../HW/src/top/ddr_tx.vhd:197:46  */
  assign n1591_o = write_request_r == write_complete_r;
  /* ../../HW/src/top/ddr_tx.vhd:197:92  */
  assign n1592_o = ~write_data_write_ena_r;
  /* ../../HW/src/top/ddr_tx.vhd:197:65  */
  assign n1593_o = n1592_o & n1591_o;
  /* ../../HW/src/top/ddr_tx.vhd:197:24  */
  assign n1594_o = n1593_o ? 1'b0 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:200:58  */
  assign n1597_o = write_addr_in[2:0];
  /* ../../HW/src/top/ddr_tx.vhd:200:43  */
  assign n1599_o = {1'b0, n1597_o};
  /* ../../HW/src/top/ddr_tx.vhd:200:104  */
  assign n1601_o = {1'b0, write_vector_in};
  /* ../../HW/src/top/ddr_tx.vhd:200:90  */
  assign n1602_o = n1599_o + n1601_o;
  /* ../../HW/src/top/ddr_tx.vhd:200:122  */
  assign n1604_o = n1602_o + 4'b0001;
  /* ../../HW/src/top/ddr_tx.vhd:200:159  */
  assign n1606_o = $unsigned(n1604_o) >= $unsigned(4'b1000);
  /* ../../HW/src/top/ddr_tx.vhd:200:23  */
  assign n1607_o = n1606_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:204:63  */
  assign n1610_o = write_addr_in[2:0];
  /* ../../HW/src/top/ddr_tx.vhd:204:48  */
  assign n1612_o = {1'b0, n1610_o};
  /* ../../HW/src/top/ddr_tx.vhd:204:109  */
  assign n1614_o = {1'b0, write_vector_in};
  /* ../../HW/src/top/ddr_tx.vhd:204:95  */
  assign n1615_o = n1612_o + n1614_o;
  /* ../../HW/src/top/ddr_tx.vhd:204:127  */
  assign n1617_o = n1615_o + 4'b0001;
  /* ../../HW/src/top/ddr_tx.vhd:204:164  */
  assign n1619_o = $unsigned(n1617_o) > $unsigned(4'b1000);
  /* ../../HW/src/top/ddr_tx.vhd:204:28  */
  assign n1620_o = n1619_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:208:53  */
  assign n1624_o = write_burstlen_in == 5'b00001;
  /* ../../HW/src/top/ddr_tx.vhd:208:95  */
  assign n1625_o = n1624_o | write_complete;
  /* ../../HW/src/top/ddr_tx.vhd:207:48  */
  assign n1626_o = n1625_o & write2;
  /* ../../HW/src/top/ddr_tx.vhd:209:34  */
  assign n1627_o = n1626_o | write_flush_r;
  /* ../../HW/src/top/ddr_tx.vhd:211:39  */
  assign n1628_o = ~hold;
  /* ../../HW/src/top/ddr_tx.vhd:210:55  */
  assign n1629_o = n1628_o & n1627_o;
  /* ../../HW/src/top/ddr_tx.vhd:207:29  */
  assign n1630_o = n1629_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:214:30  */
  assign n1632_o = ~hold;
  /* ../../HW/src/top/ddr_tx.vhd:215:43  */
  assign n1634_o = write_burstlen_in != 5'b00000;
  /* ../../HW/src/top/ddr_tx.vhd:214:35  */
  assign n1635_o = n1634_o & n1632_o;
  /* ../../HW/src/top/ddr_tx.vhd:216:38  */
  assign n1636_o = ~write_flush_r;
  /* ../../HW/src/top/ddr_tx.vhd:215:79  */
  assign n1637_o = n1636_o & n1635_o;
  /* ../../HW/src/top/ddr_tx.vhd:214:20  */
  assign n1638_o = n1637_o ? write_in : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:219:48  */
  assign n1641_o = hold | write_flush_r;
  /* ../../HW/src/top/ddr_tx.vhd:219:31  */
  assign n1642_o = n1641_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:221:60  */
  assign n1645_o = write_data_write_r[40];
  /* ../../HW/src/top/ddr_tx.vhd:221:80  */
  assign n1647_o = $unsigned(awlen_r) >= $unsigned(3'b111);
  /* ../../HW/src/top/ddr_tx.vhd:221:69  */
  assign n1648_o = n1645_o | n1647_o;
  /* ../../HW/src/top/ddr_tx.vhd:221:36  */
  assign n1649_o = n1648_o & ddr_write;
  /* ../../HW/src/top/ddr_tx.vhd:221:16  */
  assign n1650_o = n1649_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:225:17  */
  assign n1654_o = ~reset_in;
  /* ../../HW/src/top/ddr_tx.vhd:231:41  */
  assign n1657_o = awlen_r == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:231:30  */
  assign n1658_o = n1657_o & ddr_write;
  /* ../../HW/src/top/ddr_tx.vhd:232:49  */
  assign n1659_o = write_data_write_r[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:236:51  */
  assign n1662_o = write_request_r + 10'b0000000001;
  /* ../../HW/src/top/ddr_tx.vhd:238:35  */
  assign n1664_o = awlen_r + 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:237:13  */
  assign n1665_o = ddr_write ? n1664_o : awlen_r;
  /* ../../HW/src/top/ddr_tx.vhd:234:13  */
  assign n1668_o = awvalid ? 3'b000 : n1665_o;
  /* ../../HW/src/top/ddr_tx.vhd:250:21  */
  assign n1681_o = ~write_flush_r;
  /* ../../HW/src/top/ddr_tx.vhd:252:47  */
  assign n1682_o = byteenable[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:253:30  */
  assign n1683_o = {27'b0, write_burstlen_in};  //  uext
  /* ../../HW/src/top/ddr_tx.vhd:253:30  */
  assign n1685_o = n1683_o == 32'b00000000000000000000000000000001;
  /* ../../HW/src/top/ddr_tx.vhd:253:9  */
  assign n1688_o = n1685_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:260:47  */
  assign n1689_o = byteenable[7:0];
  /* ../../HW/src/top/ddr_rx.vhd:640:5  */
  assign n1691_o = {1'b1, n1689_o, write_next_addr_r};
  assign n1692_o = {n1688_o, n1682_o, wr_ddr_addr};
  /* ../../HW/src/top/ddr_tx.vhd:250:5  */
  assign n1693_o = n1681_o ? n1692_o : n1691_o;
  /* ../../HW/src/top/ddr_tx.vhd:270:129  */
  assign n1698_o = write_addr_in[31:3];
  assign n1700_o = {n1698_o, 3'b000};
  /* ../../HW/src/top/ddr_tx.vhd:277:16  */
  assign n1705_o = ~reset_in;
  /* ../../HW/src/top/ddr_tx.vhd:284:17  */
  assign n1707_o = ~hold;
  /* ../../HW/src/top/ddr_tx.vhd:289:29  */
  assign n1709_o = ~write_flush_r;
  /* ../../HW/src/top/ddr_tx.vhd:290:36  */
  assign n1711_o = write_burstlen_in == 5'b00001;
  /* ../../HW/src/top/ddr_tx.vhd:290:70  */
  assign n1712_o = write_over_complete & n1711_o;
  /* ../../HW/src/top/ddr_tx.vhd:290:16  */
  assign n1715_o = n1712_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:289:13  */
  assign n1717_o = n1709_o ? n1715_o : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:300:72  */
  assign n1720_o = wr_ddr_addr + 32'b00000000000000000000000000001000;
  /* ../../HW/src/top/ddr_tx.vhd:303:49  */
  assign n1723_o = write_complete_r + 10'b0000000001;
  /* ../../HW/src/top/ddr_tx.vhd:311:32  */
  assign n1741_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:316:35  */
  assign n1743_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:321:35  */
  assign n1745_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:321:4  */
  assign n1748_o = n1745_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/ddr_tx.vhd:321:4  */
  assign n1751_o = n1745_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/ddr_tx.vhd:321:4  */
  assign n1754_o = n1745_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/ddr_tx.vhd:316:4  */
  assign n1756_o = n1743_o ? 1'b1 : n1748_o;
  /* ../../HW/src/top/ddr_tx.vhd:316:4  */
  assign n1758_o = n1743_o ? 1'b0 : n1751_o;
  /* ../../HW/src/top/ddr_tx.vhd:316:4  */
  assign n1760_o = n1743_o ? 1'b0 : n1754_o;
  /* ../../HW/src/top/ddr_tx.vhd:311:4  */
  assign n1762_o = n1741_o ? 1'b1 : n1756_o;
  /* ../../HW/src/top/ddr_tx.vhd:311:4  */
  assign n1764_o = n1741_o ? 1'b1 : n1758_o;
  /* ../../HW/src/top/ddr_tx.vhd:311:4  */
  assign n1766_o = n1741_o ? 1'b0 : n1760_o;
  /* ../../HW/src/top/ddr_tx.vhd:334:45  */
  assign n1771_o = $unsigned(write_end_in) >= $unsigned(4'b0001);
  /* ../../HW/src/top/ddr_tx.vhd:334:26  */
  assign n1772_o = n1771_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:335:45  */
  assign n1776_o = $unsigned(write_end_in) >= $unsigned(4'b0010);
  /* ../../HW/src/top/ddr_tx.vhd:335:26  */
  assign n1777_o = n1776_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:336:45  */
  assign n1781_o = $unsigned(write_end_in) >= $unsigned(4'b0011);
  /* ../../HW/src/top/ddr_tx.vhd:336:26  */
  assign n1782_o = n1781_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:337:45  */
  assign n1786_o = $unsigned(write_end_in) >= $unsigned(4'b0100);
  /* ../../HW/src/top/ddr_tx.vhd:337:26  */
  assign n1787_o = n1786_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:338:45  */
  assign n1791_o = $unsigned(write_end_in) >= $unsigned(4'b0101);
  /* ../../HW/src/top/ddr_tx.vhd:338:26  */
  assign n1792_o = n1791_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:339:45  */
  assign n1796_o = $unsigned(write_end_in) >= $unsigned(4'b0110);
  /* ../../HW/src/top/ddr_tx.vhd:339:26  */
  assign n1797_o = n1796_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:340:45  */
  assign n1801_o = $unsigned(write_end_in) >= $unsigned(4'b0111);
  /* ../../HW/src/top/ddr_tx.vhd:340:26  */
  assign n1802_o = n1801_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:341:45  */
  assign n1806_o = $unsigned(write_end_in) >= $unsigned(4'b1000);
  /* ../../HW/src/top/ddr_tx.vhd:341:26  */
  assign n1807_o = n1806_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_tx.vhd:351:23  */
  assign n1811_o = write_addr_in[2:0];
  /* ../../HW/src/top/ddr_tx.vhd:353:103  */
  assign n1812_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:354:103  */
  assign n1813_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:355:103  */
  assign n1814_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:356:103  */
  assign n1815_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:357:103  */
  assign n1816_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:358:103  */
  assign n1817_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:359:103  */
  assign n1818_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:360:103  */
  assign n1819_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:361:100  */
  assign n1820_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:361:125  */
  assign n1821_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:361:110  */
  assign n1822_o = n1820_o | n1821_o;
  /* ../../HW/src/top/ddr_tx.vhd:362:100  */
  assign n1823_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:362:125  */
  assign n1824_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:362:110  */
  assign n1825_o = n1823_o | n1824_o;
  /* ../../HW/src/top/ddr_tx.vhd:363:100  */
  assign n1826_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:363:125  */
  assign n1827_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:363:110  */
  assign n1828_o = n1826_o | n1827_o;
  /* ../../HW/src/top/ddr_tx.vhd:364:100  */
  assign n1829_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:364:125  */
  assign n1830_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:364:110  */
  assign n1831_o = n1829_o | n1830_o;
  /* ../../HW/src/top/ddr_tx.vhd:365:100  */
  assign n1832_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:365:125  */
  assign n1833_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:365:110  */
  assign n1834_o = n1832_o | n1833_o;
  /* ../../HW/src/top/ddr_tx.vhd:366:100  */
  assign n1835_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:366:125  */
  assign n1836_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:366:110  */
  assign n1837_o = n1835_o | n1836_o;
  /* ../../HW/src/top/ddr_tx.vhd:367:100  */
  assign n1838_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:367:125  */
  assign n1839_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:367:110  */
  assign n1840_o = n1838_o | n1839_o;
  /* ../../HW/src/top/ddr_tx.vhd:368:100  */
  assign n1841_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:368:125  */
  assign n1842_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:368:110  */
  assign n1843_o = n1841_o | n1842_o;
  /* ../../HW/src/top/ddr_tx.vhd:352:9  */
  assign n1845_o = n1811_o == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:370:103  */
  assign n1846_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:371:103  */
  assign n1847_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:372:103  */
  assign n1848_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:373:103  */
  assign n1849_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:374:103  */
  assign n1850_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:375:103  */
  assign n1851_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:376:103  */
  assign n1852_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:377:100  */
  assign n1853_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:377:125  */
  assign n1854_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:377:110  */
  assign n1855_o = n1853_o | n1854_o;
  /* ../../HW/src/top/ddr_tx.vhd:378:100  */
  assign n1856_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:378:125  */
  assign n1857_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:378:110  */
  assign n1858_o = n1856_o | n1857_o;
  /* ../../HW/src/top/ddr_tx.vhd:379:100  */
  assign n1859_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:379:125  */
  assign n1860_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:379:110  */
  assign n1861_o = n1859_o | n1860_o;
  /* ../../HW/src/top/ddr_tx.vhd:380:100  */
  assign n1862_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:380:125  */
  assign n1863_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:380:110  */
  assign n1864_o = n1862_o | n1863_o;
  /* ../../HW/src/top/ddr_tx.vhd:381:100  */
  assign n1865_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:381:125  */
  assign n1866_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:381:110  */
  assign n1867_o = n1865_o | n1866_o;
  /* ../../HW/src/top/ddr_tx.vhd:382:100  */
  assign n1868_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:382:125  */
  assign n1869_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:382:110  */
  assign n1870_o = n1868_o | n1869_o;
  /* ../../HW/src/top/ddr_tx.vhd:383:100  */
  assign n1871_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:383:125  */
  assign n1872_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:383:110  */
  assign n1873_o = n1871_o | n1872_o;
  /* ../../HW/src/top/ddr_tx.vhd:384:100  */
  assign n1874_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:384:125  */
  assign n1875_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:384:110  */
  assign n1876_o = n1874_o | n1875_o;
  /* ../../HW/src/top/ddr_tx.vhd:385:103  */
  assign n1877_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:369:9  */
  assign n1879_o = n1811_o == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:387:103  */
  assign n1880_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:388:103  */
  assign n1881_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:389:103  */
  assign n1882_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:390:103  */
  assign n1883_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:391:104  */
  assign n1884_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:392:104  */
  assign n1885_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:393:101  */
  assign n1886_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:393:126  */
  assign n1887_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:393:111  */
  assign n1888_o = n1886_o | n1887_o;
  /* ../../HW/src/top/ddr_tx.vhd:394:100  */
  assign n1889_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:394:125  */
  assign n1890_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:394:110  */
  assign n1891_o = n1889_o | n1890_o;
  /* ../../HW/src/top/ddr_tx.vhd:395:100  */
  assign n1892_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:395:125  */
  assign n1893_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:395:110  */
  assign n1894_o = n1892_o | n1893_o;
  /* ../../HW/src/top/ddr_tx.vhd:396:100  */
  assign n1895_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:396:125  */
  assign n1896_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:396:110  */
  assign n1897_o = n1895_o | n1896_o;
  /* ../../HW/src/top/ddr_tx.vhd:397:100  */
  assign n1898_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:397:125  */
  assign n1899_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:397:110  */
  assign n1900_o = n1898_o | n1899_o;
  /* ../../HW/src/top/ddr_tx.vhd:398:100  */
  assign n1901_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:398:125  */
  assign n1902_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:398:110  */
  assign n1903_o = n1901_o | n1902_o;
  /* ../../HW/src/top/ddr_tx.vhd:399:100  */
  assign n1904_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:399:125  */
  assign n1905_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:399:110  */
  assign n1906_o = n1904_o | n1905_o;
  /* ../../HW/src/top/ddr_tx.vhd:400:100  */
  assign n1907_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:400:125  */
  assign n1908_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:400:110  */
  assign n1909_o = n1907_o | n1908_o;
  /* ../../HW/src/top/ddr_tx.vhd:401:103  */
  assign n1910_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:402:101  */
  assign n1911_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:386:9  */
  assign n1913_o = n1811_o == 3'b010;
  /* ../../HW/src/top/ddr_tx.vhd:404:103  */
  assign n1914_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:405:103  */
  assign n1915_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:406:103  */
  assign n1916_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:407:104  */
  assign n1917_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:408:105  */
  assign n1918_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:409:102  */
  assign n1919_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:409:127  */
  assign n1920_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:409:112  */
  assign n1921_o = n1919_o | n1920_o;
  /* ../../HW/src/top/ddr_tx.vhd:410:101  */
  assign n1922_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:410:126  */
  assign n1923_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:410:111  */
  assign n1924_o = n1922_o | n1923_o;
  /* ../../HW/src/top/ddr_tx.vhd:411:100  */
  assign n1925_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:411:125  */
  assign n1926_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:411:110  */
  assign n1927_o = n1925_o | n1926_o;
  /* ../../HW/src/top/ddr_tx.vhd:412:100  */
  assign n1928_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:412:125  */
  assign n1929_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:412:110  */
  assign n1930_o = n1928_o | n1929_o;
  /* ../../HW/src/top/ddr_tx.vhd:413:100  */
  assign n1931_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:413:125  */
  assign n1932_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:413:110  */
  assign n1933_o = n1931_o | n1932_o;
  /* ../../HW/src/top/ddr_tx.vhd:414:100  */
  assign n1934_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:414:125  */
  assign n1935_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:414:110  */
  assign n1936_o = n1934_o | n1935_o;
  /* ../../HW/src/top/ddr_tx.vhd:415:100  */
  assign n1937_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:415:125  */
  assign n1938_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:415:110  */
  assign n1939_o = n1937_o | n1938_o;
  /* ../../HW/src/top/ddr_tx.vhd:416:100  */
  assign n1940_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:416:125  */
  assign n1941_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:416:110  */
  assign n1942_o = n1940_o | n1941_o;
  /* ../../HW/src/top/ddr_tx.vhd:417:103  */
  assign n1943_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:418:101  */
  assign n1944_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:419:101  */
  assign n1945_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:403:9  */
  assign n1947_o = n1811_o == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:421:103  */
  assign n1948_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:422:103  */
  assign n1949_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:423:104  */
  assign n1950_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:424:105  */
  assign n1951_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:425:102  */
  assign n1952_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:425:127  */
  assign n1953_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:425:112  */
  assign n1954_o = n1952_o | n1953_o;
  /* ../../HW/src/top/ddr_tx.vhd:426:102  */
  assign n1955_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:426:127  */
  assign n1956_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:426:112  */
  assign n1957_o = n1955_o | n1956_o;
  /* ../../HW/src/top/ddr_tx.vhd:427:101  */
  assign n1958_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:427:126  */
  assign n1959_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:427:111  */
  assign n1960_o = n1958_o | n1959_o;
  /* ../../HW/src/top/ddr_tx.vhd:428:100  */
  assign n1961_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:428:125  */
  assign n1962_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:428:110  */
  assign n1963_o = n1961_o | n1962_o;
  /* ../../HW/src/top/ddr_tx.vhd:429:100  */
  assign n1964_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:429:125  */
  assign n1965_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:429:110  */
  assign n1966_o = n1964_o | n1965_o;
  /* ../../HW/src/top/ddr_tx.vhd:430:100  */
  assign n1967_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:430:125  */
  assign n1968_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:430:110  */
  assign n1969_o = n1967_o | n1968_o;
  /* ../../HW/src/top/ddr_tx.vhd:431:100  */
  assign n1970_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:431:125  */
  assign n1971_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:431:110  */
  assign n1972_o = n1970_o | n1971_o;
  /* ../../HW/src/top/ddr_tx.vhd:432:100  */
  assign n1973_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:432:125  */
  assign n1974_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:432:110  */
  assign n1975_o = n1973_o | n1974_o;
  /* ../../HW/src/top/ddr_tx.vhd:433:103  */
  assign n1976_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:434:101  */
  assign n1977_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:435:101  */
  assign n1978_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:436:101  */
  assign n1979_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:420:9  */
  assign n1981_o = n1811_o == 3'b100;
  /* ../../HW/src/top/ddr_tx.vhd:438:103  */
  assign n1982_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:439:104  */
  assign n1983_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:440:105  */
  assign n1984_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:441:102  */
  assign n1985_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:441:127  */
  assign n1986_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:441:112  */
  assign n1987_o = n1985_o | n1986_o;
  /* ../../HW/src/top/ddr_tx.vhd:442:102  */
  assign n1988_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:442:127  */
  assign n1989_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:442:112  */
  assign n1990_o = n1988_o | n1989_o;
  /* ../../HW/src/top/ddr_tx.vhd:443:102  */
  assign n1991_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:443:127  */
  assign n1992_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:443:112  */
  assign n1993_o = n1991_o | n1992_o;
  /* ../../HW/src/top/ddr_tx.vhd:444:101  */
  assign n1994_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:444:126  */
  assign n1995_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:444:111  */
  assign n1996_o = n1994_o | n1995_o;
  /* ../../HW/src/top/ddr_tx.vhd:445:100  */
  assign n1997_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:445:125  */
  assign n1998_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:445:110  */
  assign n1999_o = n1997_o | n1998_o;
  /* ../../HW/src/top/ddr_tx.vhd:446:100  */
  assign n2000_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:446:125  */
  assign n2001_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:446:110  */
  assign n2002_o = n2000_o | n2001_o;
  /* ../../HW/src/top/ddr_tx.vhd:447:100  */
  assign n2003_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:447:125  */
  assign n2004_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:447:110  */
  assign n2005_o = n2003_o | n2004_o;
  /* ../../HW/src/top/ddr_tx.vhd:448:100  */
  assign n2006_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:448:125  */
  assign n2007_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:448:110  */
  assign n2008_o = n2006_o | n2007_o;
  /* ../../HW/src/top/ddr_tx.vhd:449:103  */
  assign n2009_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:450:101  */
  assign n2010_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:451:101  */
  assign n2011_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:452:101  */
  assign n2012_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:453:101  */
  assign n2013_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:437:9  */
  assign n2015_o = n1811_o == 3'b101;
  /* ../../HW/src/top/ddr_tx.vhd:455:104  */
  assign n2016_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:456:105  */
  assign n2017_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:457:102  */
  assign n2018_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:457:127  */
  assign n2019_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:457:112  */
  assign n2020_o = n2018_o | n2019_o;
  /* ../../HW/src/top/ddr_tx.vhd:458:102  */
  assign n2021_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:458:127  */
  assign n2022_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:458:112  */
  assign n2023_o = n2021_o | n2022_o;
  /* ../../HW/src/top/ddr_tx.vhd:459:102  */
  assign n2024_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:459:127  */
  assign n2025_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:459:112  */
  assign n2026_o = n2024_o | n2025_o;
  /* ../../HW/src/top/ddr_tx.vhd:460:102  */
  assign n2027_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:460:127  */
  assign n2028_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:460:112  */
  assign n2029_o = n2027_o | n2028_o;
  /* ../../HW/src/top/ddr_tx.vhd:461:101  */
  assign n2030_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:461:126  */
  assign n2031_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:461:111  */
  assign n2032_o = n2030_o | n2031_o;
  /* ../../HW/src/top/ddr_tx.vhd:462:100  */
  assign n2033_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:462:125  */
  assign n2034_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:462:110  */
  assign n2035_o = n2033_o | n2034_o;
  /* ../../HW/src/top/ddr_tx.vhd:463:100  */
  assign n2036_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:463:125  */
  assign n2037_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:463:110  */
  assign n2038_o = n2036_o | n2037_o;
  /* ../../HW/src/top/ddr_tx.vhd:464:100  */
  assign n2039_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:464:125  */
  assign n2040_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:464:110  */
  assign n2041_o = n2039_o | n2040_o;
  /* ../../HW/src/top/ddr_tx.vhd:465:103  */
  assign n2042_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:466:101  */
  assign n2043_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:467:101  */
  assign n2044_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:468:101  */
  assign n2045_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:469:101  */
  assign n2046_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:470:101  */
  assign n2047_o = byteenable_r[0];
  /* ../../HW/src/top/ddr_tx.vhd:454:9  */
  assign n2049_o = n1811_o == 3'b110;
  /* ../../HW/src/top/ddr_tx.vhd:472:105  */
  assign n2050_o = byteenable_r[15];
  /* ../../HW/src/top/ddr_tx.vhd:473:102  */
  assign n2051_o = w_mask8 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:473:127  */
  assign n2052_o = byteenable_r[14];
  /* ../../HW/src/top/ddr_tx.vhd:473:112  */
  assign n2053_o = n2051_o | n2052_o;
  /* ../../HW/src/top/ddr_tx.vhd:474:102  */
  assign n2054_o = w_mask7 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:474:127  */
  assign n2055_o = byteenable_r[13];
  /* ../../HW/src/top/ddr_tx.vhd:474:112  */
  assign n2056_o = n2054_o | n2055_o;
  /* ../../HW/src/top/ddr_tx.vhd:475:102  */
  assign n2057_o = w_mask6 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:475:127  */
  assign n2058_o = byteenable_r[12];
  /* ../../HW/src/top/ddr_tx.vhd:475:112  */
  assign n2059_o = n2057_o | n2058_o;
  /* ../../HW/src/top/ddr_tx.vhd:476:102  */
  assign n2060_o = w_mask5 & w_x8;
  /* ../../HW/src/top/ddr_tx.vhd:476:127  */
  assign n2061_o = byteenable_r[11];
  /* ../../HW/src/top/ddr_tx.vhd:476:112  */
  assign n2062_o = n2060_o | n2061_o;
  /* ../../HW/src/top/ddr_tx.vhd:477:102  */
  assign n2063_o = w_mask4 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:477:127  */
  assign n2064_o = byteenable_r[10];
  /* ../../HW/src/top/ddr_tx.vhd:477:112  */
  assign n2065_o = n2063_o | n2064_o;
  /* ../../HW/src/top/ddr_tx.vhd:478:101  */
  assign n2066_o = w_mask3 & w_x4;
  /* ../../HW/src/top/ddr_tx.vhd:478:126  */
  assign n2067_o = byteenable_r[9];
  /* ../../HW/src/top/ddr_tx.vhd:478:111  */
  assign n2068_o = n2066_o | n2067_o;
  /* ../../HW/src/top/ddr_tx.vhd:479:100  */
  assign n2069_o = w_mask2 & w_x2;
  /* ../../HW/src/top/ddr_tx.vhd:479:125  */
  assign n2070_o = byteenable_r[8];
  /* ../../HW/src/top/ddr_tx.vhd:479:110  */
  assign n2071_o = n2069_o | n2070_o;
  /* ../../HW/src/top/ddr_tx.vhd:480:100  */
  assign n2072_o = w_mask1 & w_x1;
  /* ../../HW/src/top/ddr_tx.vhd:480:125  */
  assign n2073_o = byteenable_r[7];
  /* ../../HW/src/top/ddr_tx.vhd:480:110  */
  assign n2074_o = n2072_o | n2073_o;
  /* ../../HW/src/top/ddr_tx.vhd:481:103  */
  assign n2075_o = byteenable_r[6];
  /* ../../HW/src/top/ddr_tx.vhd:482:101  */
  assign n2076_o = byteenable_r[5];
  /* ../../HW/src/top/ddr_tx.vhd:483:101  */
  assign n2077_o = byteenable_r[4];
  /* ../../HW/src/top/ddr_tx.vhd:484:101  */
  assign n2078_o = byteenable_r[3];
  /* ../../HW/src/top/ddr_tx.vhd:485:101  */
  assign n2079_o = byteenable_r[2];
  /* ../../HW/src/top/ddr_tx.vhd:486:101  */
  assign n2080_o = byteenable_r[1];
  /* ../../HW/src/top/ddr_tx.vhd:487:102  */
  assign n2081_o = byteenable_r[0];
  assign n2082_o = {n2049_o, n2015_o, n1981_o, n1947_o, n1913_o, n1879_o, n1845_o};
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2083_o = n2047_o;
      7'b0100000: n2083_o = n2013_o;
      7'b0010000: n2083_o = n1979_o;
      7'b0001000: n2083_o = n1945_o;
      7'b0000100: n2083_o = n1911_o;
      7'b0000010: n2083_o = n1877_o;
      7'b0000001: n2083_o = n1843_o;
      default: n2083_o = n2081_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2084_o = n2046_o;
      7'b0100000: n2084_o = n2012_o;
      7'b0010000: n2084_o = n1978_o;
      7'b0001000: n2084_o = n1944_o;
      7'b0000100: n2084_o = n1910_o;
      7'b0000010: n2084_o = n1876_o;
      7'b0000001: n2084_o = n1840_o;
      default: n2084_o = n2080_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2085_o = n2045_o;
      7'b0100000: n2085_o = n2011_o;
      7'b0010000: n2085_o = n1977_o;
      7'b0001000: n2085_o = n1943_o;
      7'b0000100: n2085_o = n1909_o;
      7'b0000010: n2085_o = n1873_o;
      7'b0000001: n2085_o = n1837_o;
      default: n2085_o = n2079_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2086_o = n2044_o;
      7'b0100000: n2086_o = n2010_o;
      7'b0010000: n2086_o = n1976_o;
      7'b0001000: n2086_o = n1942_o;
      7'b0000100: n2086_o = n1906_o;
      7'b0000010: n2086_o = n1870_o;
      7'b0000001: n2086_o = n1834_o;
      default: n2086_o = n2078_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2087_o = n2043_o;
      7'b0100000: n2087_o = n2009_o;
      7'b0010000: n2087_o = n1975_o;
      7'b0001000: n2087_o = n1939_o;
      7'b0000100: n2087_o = n1903_o;
      7'b0000010: n2087_o = n1867_o;
      7'b0000001: n2087_o = n1831_o;
      default: n2087_o = n2077_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2088_o = n2042_o;
      7'b0100000: n2088_o = n2008_o;
      7'b0010000: n2088_o = n1972_o;
      7'b0001000: n2088_o = n1936_o;
      7'b0000100: n2088_o = n1900_o;
      7'b0000010: n2088_o = n1864_o;
      7'b0000001: n2088_o = n1828_o;
      default: n2088_o = n2076_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2089_o = n2041_o;
      7'b0100000: n2089_o = n2005_o;
      7'b0010000: n2089_o = n1969_o;
      7'b0001000: n2089_o = n1933_o;
      7'b0000100: n2089_o = n1897_o;
      7'b0000010: n2089_o = n1861_o;
      7'b0000001: n2089_o = n1825_o;
      default: n2089_o = n2075_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2090_o = n2038_o;
      7'b0100000: n2090_o = n2002_o;
      7'b0010000: n2090_o = n1966_o;
      7'b0001000: n2090_o = n1930_o;
      7'b0000100: n2090_o = n1894_o;
      7'b0000010: n2090_o = n1858_o;
      7'b0000001: n2090_o = n1822_o;
      default: n2090_o = n2074_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2091_o = n2035_o;
      7'b0100000: n2091_o = n1999_o;
      7'b0010000: n2091_o = n1963_o;
      7'b0001000: n2091_o = n1927_o;
      7'b0000100: n2091_o = n1891_o;
      7'b0000010: n2091_o = n1855_o;
      7'b0000001: n2091_o = n1819_o;
      default: n2091_o = n2071_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2092_o = n2032_o;
      7'b0100000: n2092_o = n1996_o;
      7'b0010000: n2092_o = n1960_o;
      7'b0001000: n2092_o = n1924_o;
      7'b0000100: n2092_o = n1888_o;
      7'b0000010: n2092_o = n1852_o;
      7'b0000001: n2092_o = n1818_o;
      default: n2092_o = n2068_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2093_o = n2029_o;
      7'b0100000: n2093_o = n1993_o;
      7'b0010000: n2093_o = n1957_o;
      7'b0001000: n2093_o = n1921_o;
      7'b0000100: n2093_o = n1885_o;
      7'b0000010: n2093_o = n1851_o;
      7'b0000001: n2093_o = n1817_o;
      default: n2093_o = n2065_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2094_o = n2026_o;
      7'b0100000: n2094_o = n1990_o;
      7'b0010000: n2094_o = n1954_o;
      7'b0001000: n2094_o = n1918_o;
      7'b0000100: n2094_o = n1884_o;
      7'b0000010: n2094_o = n1850_o;
      7'b0000001: n2094_o = n1816_o;
      default: n2094_o = n2062_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2095_o = n2023_o;
      7'b0100000: n2095_o = n1987_o;
      7'b0010000: n2095_o = n1951_o;
      7'b0001000: n2095_o = n1917_o;
      7'b0000100: n2095_o = n1883_o;
      7'b0000010: n2095_o = n1849_o;
      7'b0000001: n2095_o = n1815_o;
      default: n2095_o = n2059_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2096_o = n2020_o;
      7'b0100000: n2096_o = n1984_o;
      7'b0010000: n2096_o = n1950_o;
      7'b0001000: n2096_o = n1916_o;
      7'b0000100: n2096_o = n1882_o;
      7'b0000010: n2096_o = n1848_o;
      7'b0000001: n2096_o = n1814_o;
      default: n2096_o = n2056_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2097_o = n2017_o;
      7'b0100000: n2097_o = n1983_o;
      7'b0010000: n2097_o = n1949_o;
      7'b0001000: n2097_o = n1915_o;
      7'b0000100: n2097_o = n1881_o;
      7'b0000010: n2097_o = n1847_o;
      7'b0000001: n2097_o = n1813_o;
      default: n2097_o = n2053_o;
    endcase
  /* ../../HW/src/top/ddr_tx.vhd:351:5  */
  always @*
    case (n2082_o)
      7'b1000000: n2098_o = n2016_o;
      7'b0100000: n2098_o = n1982_o;
      7'b0010000: n2098_o = n1948_o;
      7'b0001000: n2098_o = n1914_o;
      7'b0000100: n2098_o = n1880_o;
      7'b0000010: n2098_o = n1846_o;
      7'b0000001: n2098_o = n1812_o;
      default: n2098_o = n2050_o;
    endcase
  assign n2099_o = {n2098_o, n2097_o, n2096_o, n2095_o, n2094_o, n2093_o, n2092_o, n2091_o, n2090_o, n2089_o, n2088_o, n2087_o, n2086_o, n2085_o, n2084_o, n2083_o};
  /* ../../HW/src/top/ddr_tx.vhd:350:1  */
  assign n2100_o = write2 ? n2099_o : byteenable_r;
  /* ../../HW/src/top/ddr_tx.vhd:498:23  */
  assign n2104_o = write_addr_in[2:0];
  /* ../../HW/src/top/ddr_tx.vhd:500:41  */
  assign n2106_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:501:115  */
  assign n2107_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:502:44  */
  assign n2109_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:503:115  */
  assign n2110_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:504:44  */
  assign n2112_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:505:115  */
  assign n2113_o = write_data_in[7:0];
  assign n2114_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:504:13  */
  assign n2115_o = n2112_o ? n2113_o : n2114_o;
  assign n2116_o = write_data_in[63:8];
  assign n2117_o = write_data_r[63:8];
  /* ../../HW/src/top/ddr_tx.vhd:504:13  */
  assign n2118_o = n2112_o ? n2117_o : n2116_o;
  assign n2119_o = {n2118_o, n2115_o};
  assign n2120_o = n2119_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:502:13  */
  assign n2121_o = n2109_o ? n2110_o : n2120_o;
  assign n2122_o = n2119_o[63:16];
  assign n2123_o = write_data_r[63:16];
  /* ../../HW/src/top/ddr_tx.vhd:502:13  */
  assign n2124_o = n2109_o ? n2123_o : n2122_o;
  assign n2125_o = {n2124_o, n2121_o};
  assign n2126_o = n2125_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:500:13  */
  assign n2127_o = n2106_o ? n2107_o : n2126_o;
  assign n2128_o = n2125_o[63:32];
  assign n2129_o = write_data_r[63:32];
  /* ../../HW/src/top/ddr_tx.vhd:500:13  */
  assign n2130_o = n2106_o ? n2129_o : n2128_o;
  /* ../../HW/src/top/ddr_tx.vhd:499:9  */
  assign n2132_o = n2104_o == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:510:41  */
  assign n2134_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:511:115  */
  assign n2135_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:512:44  */
  assign n2137_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:513:115  */
  assign n2138_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:514:44  */
  assign n2140_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:515:115  */
  assign n2141_o = write_data_in[7:0];
  assign n2142_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:514:13  */
  assign n2143_o = n2140_o ? n2141_o : n2142_o;
  assign n2144_o = write_data_in[63:8];
  assign n2145_o = write_data_r[71:16];
  /* ../../HW/src/top/ddr_tx.vhd:514:13  */
  assign n2146_o = n2140_o ? n2145_o : n2144_o;
  assign n2147_o = {n2146_o, n2143_o};
  assign n2148_o = n2147_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:512:13  */
  assign n2149_o = n2137_o ? n2138_o : n2148_o;
  assign n2150_o = n2147_o[63:16];
  assign n2151_o = write_data_r[71:24];
  /* ../../HW/src/top/ddr_tx.vhd:512:13  */
  assign n2152_o = n2137_o ? n2151_o : n2150_o;
  assign n2153_o = {n2152_o, n2149_o};
  assign n2154_o = n2153_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:510:13  */
  assign n2155_o = n2134_o ? n2135_o : n2154_o;
  assign n2156_o = n2153_o[63:32];
  assign n2157_o = write_data_r[71:40];
  /* ../../HW/src/top/ddr_tx.vhd:510:13  */
  assign n2158_o = n2134_o ? n2157_o : n2156_o;
  /* ../../HW/src/top/ddr_tx.vhd:509:9  */
  assign n2160_o = n2104_o == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:520:41  */
  assign n2162_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:521:115  */
  assign n2163_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:522:44  */
  assign n2165_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:523:115  */
  assign n2166_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:524:44  */
  assign n2168_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:525:114  */
  assign n2169_o = write_data_in[7:0];
  assign n2170_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:524:13  */
  assign n2171_o = n2168_o ? n2169_o : n2170_o;
  assign n2172_o = write_data_in[63:8];
  assign n2173_o = write_data_r[79:24];
  /* ../../HW/src/top/ddr_tx.vhd:524:13  */
  assign n2174_o = n2168_o ? n2173_o : n2172_o;
  assign n2175_o = {n2174_o, n2171_o};
  assign n2176_o = n2175_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:522:13  */
  assign n2177_o = n2165_o ? n2166_o : n2176_o;
  assign n2178_o = n2175_o[63:16];
  assign n2179_o = write_data_r[79:32];
  /* ../../HW/src/top/ddr_tx.vhd:522:13  */
  assign n2180_o = n2165_o ? n2179_o : n2178_o;
  assign n2181_o = {n2180_o, n2177_o};
  assign n2182_o = n2181_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:520:13  */
  assign n2183_o = n2162_o ? n2163_o : n2182_o;
  assign n2184_o = n2181_o[63:32];
  assign n2185_o = write_data_r[79:48];
  /* ../../HW/src/top/ddr_tx.vhd:520:13  */
  assign n2186_o = n2162_o ? n2185_o : n2184_o;
  /* ../../HW/src/top/ddr_tx.vhd:519:9  */
  assign n2188_o = n2104_o == 3'b010;
  /* ../../HW/src/top/ddr_tx.vhd:530:41  */
  assign n2190_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:531:115  */
  assign n2191_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:532:44  */
  assign n2193_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:533:115  */
  assign n2194_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:534:44  */
  assign n2196_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:535:114  */
  assign n2197_o = write_data_in[7:0];
  assign n2198_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:534:13  */
  assign n2199_o = n2196_o ? n2197_o : n2198_o;
  assign n2200_o = write_data_in[63:8];
  assign n2201_o = write_data_r[87:32];
  /* ../../HW/src/top/ddr_tx.vhd:534:13  */
  assign n2202_o = n2196_o ? n2201_o : n2200_o;
  assign n2203_o = {n2202_o, n2199_o};
  assign n2204_o = n2203_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:532:13  */
  assign n2205_o = n2193_o ? n2194_o : n2204_o;
  assign n2206_o = n2203_o[63:16];
  assign n2207_o = write_data_r[87:40];
  /* ../../HW/src/top/ddr_tx.vhd:532:13  */
  assign n2208_o = n2193_o ? n2207_o : n2206_o;
  assign n2209_o = {n2208_o, n2205_o};
  assign n2210_o = n2209_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:530:13  */
  assign n2211_o = n2190_o ? n2191_o : n2210_o;
  assign n2212_o = n2209_o[63:32];
  assign n2213_o = write_data_r[87:56];
  /* ../../HW/src/top/ddr_tx.vhd:530:13  */
  assign n2214_o = n2190_o ? n2213_o : n2212_o;
  /* ../../HW/src/top/ddr_tx.vhd:529:9  */
  assign n2216_o = n2104_o == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:540:41  */
  assign n2218_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:541:115  */
  assign n2219_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:542:44  */
  assign n2221_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:543:115  */
  assign n2222_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:544:44  */
  assign n2224_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:545:114  */
  assign n2225_o = write_data_in[7:0];
  assign n2226_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:544:13  */
  assign n2227_o = n2224_o ? n2225_o : n2226_o;
  assign n2228_o = write_data_in[63:8];
  assign n2229_o = write_data_r[95:40];
  /* ../../HW/src/top/ddr_tx.vhd:544:13  */
  assign n2230_o = n2224_o ? n2229_o : n2228_o;
  assign n2231_o = {n2230_o, n2227_o};
  assign n2232_o = n2231_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:542:13  */
  assign n2233_o = n2221_o ? n2222_o : n2232_o;
  assign n2234_o = n2231_o[63:16];
  assign n2235_o = write_data_r[95:48];
  /* ../../HW/src/top/ddr_tx.vhd:542:13  */
  assign n2236_o = n2221_o ? n2235_o : n2234_o;
  assign n2237_o = {n2236_o, n2233_o};
  assign n2238_o = n2237_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:540:13  */
  assign n2239_o = n2218_o ? n2219_o : n2238_o;
  assign n2240_o = n2237_o[63:32];
  assign n2241_o = write_data_r[95:64];
  /* ../../HW/src/top/ddr_tx.vhd:540:13  */
  assign n2242_o = n2218_o ? n2241_o : n2240_o;
  /* ../../HW/src/top/ddr_tx.vhd:539:9  */
  assign n2244_o = n2104_o == 3'b100;
  /* ../../HW/src/top/ddr_tx.vhd:550:41  */
  assign n2246_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:551:115  */
  assign n2247_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:552:44  */
  assign n2249_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:553:115  */
  assign n2250_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:554:44  */
  assign n2252_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:555:114  */
  assign n2253_o = write_data_in[7:0];
  assign n2254_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:554:13  */
  assign n2255_o = n2252_o ? n2253_o : n2254_o;
  assign n2256_o = write_data_in[63:8];
  assign n2257_o = write_data_r[103:48];
  /* ../../HW/src/top/ddr_tx.vhd:554:13  */
  assign n2258_o = n2252_o ? n2257_o : n2256_o;
  assign n2259_o = {n2258_o, n2255_o};
  assign n2260_o = n2259_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:552:13  */
  assign n2261_o = n2249_o ? n2250_o : n2260_o;
  assign n2262_o = n2259_o[63:16];
  assign n2263_o = write_data_r[103:56];
  /* ../../HW/src/top/ddr_tx.vhd:552:13  */
  assign n2264_o = n2249_o ? n2263_o : n2262_o;
  assign n2265_o = {n2264_o, n2261_o};
  assign n2266_o = n2265_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:550:13  */
  assign n2267_o = n2246_o ? n2247_o : n2266_o;
  assign n2268_o = n2265_o[63:32];
  assign n2269_o = write_data_r[103:72];
  /* ../../HW/src/top/ddr_tx.vhd:550:13  */
  assign n2270_o = n2246_o ? n2269_o : n2268_o;
  /* ../../HW/src/top/ddr_tx.vhd:549:9  */
  assign n2272_o = n2104_o == 3'b101;
  /* ../../HW/src/top/ddr_tx.vhd:560:41  */
  assign n2274_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:561:115  */
  assign n2275_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:562:44  */
  assign n2277_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:563:115  */
  assign n2278_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:564:44  */
  assign n2280_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:565:114  */
  assign n2281_o = write_data_in[7:0];
  assign n2282_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:564:13  */
  assign n2283_o = n2280_o ? n2281_o : n2282_o;
  assign n2284_o = write_data_in[63:8];
  assign n2285_o = write_data_r[111:56];
  /* ../../HW/src/top/ddr_tx.vhd:564:13  */
  assign n2286_o = n2280_o ? n2285_o : n2284_o;
  assign n2287_o = {n2286_o, n2283_o};
  assign n2288_o = n2287_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:562:13  */
  assign n2289_o = n2277_o ? n2278_o : n2288_o;
  assign n2290_o = n2287_o[63:16];
  assign n2291_o = write_data_r[111:64];
  /* ../../HW/src/top/ddr_tx.vhd:562:13  */
  assign n2292_o = n2277_o ? n2291_o : n2290_o;
  assign n2293_o = {n2292_o, n2289_o};
  assign n2294_o = n2293_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:560:13  */
  assign n2295_o = n2274_o ? n2275_o : n2294_o;
  assign n2296_o = n2293_o[63:32];
  assign n2297_o = write_data_r[111:80];
  /* ../../HW/src/top/ddr_tx.vhd:560:13  */
  assign n2298_o = n2274_o ? n2297_o : n2296_o;
  /* ../../HW/src/top/ddr_tx.vhd:559:9  */
  assign n2300_o = n2104_o == 3'b110;
  /* ../../HW/src/top/ddr_tx.vhd:570:41  */
  assign n2302_o = write_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_tx.vhd:571:115  */
  assign n2303_o = write_data_in[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:572:44  */
  assign n2305_o = write_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_tx.vhd:573:115  */
  assign n2306_o = write_data_in[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:574:44  */
  assign n2308_o = write_vector_in == 3'b000;
  /* ../../HW/src/top/ddr_tx.vhd:575:114  */
  assign n2309_o = write_data_in[7:0];
  assign n2310_o = write_data_in[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:574:13  */
  assign n2311_o = n2308_o ? n2309_o : n2310_o;
  assign n2312_o = write_data_in[63:8];
  assign n2313_o = write_data_r[119:64];
  /* ../../HW/src/top/ddr_tx.vhd:574:13  */
  assign n2314_o = n2308_o ? n2313_o : n2312_o;
  assign n2315_o = {n2314_o, n2311_o};
  assign n2316_o = n2315_o[15:0];
  /* ../../HW/src/top/ddr_tx.vhd:572:13  */
  assign n2317_o = n2305_o ? n2306_o : n2316_o;
  assign n2318_o = n2315_o[63:16];
  assign n2319_o = write_data_r[119:72];
  /* ../../HW/src/top/ddr_tx.vhd:572:13  */
  assign n2320_o = n2305_o ? n2319_o : n2318_o;
  assign n2321_o = {n2320_o, n2317_o};
  assign n2322_o = n2321_o[31:0];
  /* ../../HW/src/top/ddr_tx.vhd:570:13  */
  assign n2323_o = n2302_o ? n2303_o : n2322_o;
  assign n2324_o = n2321_o[63:32];
  assign n2325_o = write_data_r[119:88];
  /* ../../HW/src/top/ddr_tx.vhd:570:13  */
  assign n2326_o = n2302_o ? n2325_o : n2324_o;
  assign n2327_o = {n2300_o, n2272_o, n2244_o, n2216_o, n2188_o, n2160_o, n2132_o};
  assign n2328_o = n2127_o[7:0];
  assign n2329_o = write_data_r[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2330_o = n2329_o;
      7'b0100000: n2330_o = n2329_o;
      7'b0010000: n2330_o = n2329_o;
      7'b0001000: n2330_o = n2329_o;
      7'b0000100: n2330_o = n2329_o;
      7'b0000010: n2330_o = n2329_o;
      7'b0000001: n2330_o = n2328_o;
      default: n2330_o = n2329_o;
    endcase
  assign n2331_o = n2127_o[15:8];
  assign n2332_o = n2155_o[7:0];
  assign n2333_o = write_data_r[15:8];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2334_o = n2333_o;
      7'b0100000: n2334_o = n2333_o;
      7'b0010000: n2334_o = n2333_o;
      7'b0001000: n2334_o = n2333_o;
      7'b0000100: n2334_o = n2333_o;
      7'b0000010: n2334_o = n2332_o;
      7'b0000001: n2334_o = n2331_o;
      default: n2334_o = n2333_o;
    endcase
  assign n2335_o = n2127_o[23:16];
  assign n2336_o = n2155_o[15:8];
  assign n2337_o = n2183_o[7:0];
  assign n2338_o = write_data_r[23:16];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2339_o = n2338_o;
      7'b0100000: n2339_o = n2338_o;
      7'b0010000: n2339_o = n2338_o;
      7'b0001000: n2339_o = n2338_o;
      7'b0000100: n2339_o = n2337_o;
      7'b0000010: n2339_o = n2336_o;
      7'b0000001: n2339_o = n2335_o;
      default: n2339_o = n2338_o;
    endcase
  assign n2340_o = n2127_o[31:24];
  assign n2341_o = n2155_o[23:16];
  assign n2342_o = n2183_o[15:8];
  assign n2343_o = n2211_o[7:0];
  assign n2344_o = write_data_r[31:24];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2345_o = n2344_o;
      7'b0100000: n2345_o = n2344_o;
      7'b0010000: n2345_o = n2344_o;
      7'b0001000: n2345_o = n2343_o;
      7'b0000100: n2345_o = n2342_o;
      7'b0000010: n2345_o = n2341_o;
      7'b0000001: n2345_o = n2340_o;
      default: n2345_o = n2344_o;
    endcase
  assign n2346_o = n2130_o[7:0];
  assign n2347_o = n2155_o[31:24];
  assign n2348_o = n2183_o[23:16];
  assign n2349_o = n2211_o[15:8];
  assign n2350_o = n2239_o[7:0];
  assign n2351_o = write_data_r[39:32];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2352_o = n2351_o;
      7'b0100000: n2352_o = n2351_o;
      7'b0010000: n2352_o = n2350_o;
      7'b0001000: n2352_o = n2349_o;
      7'b0000100: n2352_o = n2348_o;
      7'b0000010: n2352_o = n2347_o;
      7'b0000001: n2352_o = n2346_o;
      default: n2352_o = n2351_o;
    endcase
  assign n2353_o = n2130_o[15:8];
  assign n2354_o = n2158_o[7:0];
  assign n2355_o = n2183_o[31:24];
  assign n2356_o = n2211_o[23:16];
  assign n2357_o = n2239_o[15:8];
  assign n2358_o = n2267_o[7:0];
  assign n2359_o = write_data_r[47:40];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2360_o = n2359_o;
      7'b0100000: n2360_o = n2358_o;
      7'b0010000: n2360_o = n2357_o;
      7'b0001000: n2360_o = n2356_o;
      7'b0000100: n2360_o = n2355_o;
      7'b0000010: n2360_o = n2354_o;
      7'b0000001: n2360_o = n2353_o;
      default: n2360_o = n2359_o;
    endcase
  assign n2361_o = n2130_o[23:16];
  assign n2362_o = n2158_o[15:8];
  assign n2363_o = n2186_o[7:0];
  assign n2364_o = n2211_o[31:24];
  assign n2365_o = n2239_o[23:16];
  assign n2366_o = n2267_o[15:8];
  assign n2367_o = n2295_o[7:0];
  assign n2368_o = write_data_r[55:48];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2369_o = n2367_o;
      7'b0100000: n2369_o = n2366_o;
      7'b0010000: n2369_o = n2365_o;
      7'b0001000: n2369_o = n2364_o;
      7'b0000100: n2369_o = n2363_o;
      7'b0000010: n2369_o = n2362_o;
      7'b0000001: n2369_o = n2361_o;
      default: n2369_o = n2368_o;
    endcase
  assign n2370_o = n2130_o[31:24];
  assign n2371_o = n2158_o[23:16];
  assign n2372_o = n2186_o[15:8];
  assign n2373_o = n2214_o[7:0];
  assign n2374_o = n2239_o[31:24];
  assign n2375_o = n2267_o[23:16];
  assign n2376_o = n2295_o[15:8];
  assign n2377_o = n2323_o[7:0];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2378_o = n2376_o;
      7'b0100000: n2378_o = n2375_o;
      7'b0010000: n2378_o = n2374_o;
      7'b0001000: n2378_o = n2373_o;
      7'b0000100: n2378_o = n2372_o;
      7'b0000010: n2378_o = n2371_o;
      7'b0000001: n2378_o = n2370_o;
      default: n2378_o = n2377_o;
    endcase
  assign n2379_o = n2158_o[31:24];
  assign n2380_o = n2186_o[23:16];
  assign n2381_o = n2214_o[15:8];
  assign n2382_o = n2242_o[7:0];
  assign n2383_o = n2267_o[31:24];
  assign n2384_o = n2295_o[23:16];
  assign n2385_o = n2323_o[15:8];
  assign n2386_o = write_data_r[71:64];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2387_o = n2384_o;
      7'b0100000: n2387_o = n2383_o;
      7'b0010000: n2387_o = n2382_o;
      7'b0001000: n2387_o = n2381_o;
      7'b0000100: n2387_o = n2380_o;
      7'b0000010: n2387_o = n2379_o;
      7'b0000001: n2387_o = n2386_o;
      default: n2387_o = n2385_o;
    endcase
  assign n2388_o = n2186_o[31:24];
  assign n2389_o = n2214_o[23:16];
  assign n2390_o = n2242_o[15:8];
  assign n2391_o = n2270_o[7:0];
  assign n2392_o = n2295_o[31:24];
  assign n2393_o = n2323_o[23:16];
  assign n2394_o = write_data_r[79:72];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2395_o = n2392_o;
      7'b0100000: n2395_o = n2391_o;
      7'b0010000: n2395_o = n2390_o;
      7'b0001000: n2395_o = n2389_o;
      7'b0000100: n2395_o = n2388_o;
      7'b0000010: n2395_o = n2394_o;
      7'b0000001: n2395_o = n2394_o;
      default: n2395_o = n2393_o;
    endcase
  assign n2396_o = n2214_o[31:24];
  assign n2397_o = n2242_o[23:16];
  assign n2398_o = n2270_o[15:8];
  assign n2399_o = n2298_o[7:0];
  assign n2400_o = n2323_o[31:24];
  assign n2401_o = write_data_r[87:80];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2402_o = n2399_o;
      7'b0100000: n2402_o = n2398_o;
      7'b0010000: n2402_o = n2397_o;
      7'b0001000: n2402_o = n2396_o;
      7'b0000100: n2402_o = n2401_o;
      7'b0000010: n2402_o = n2401_o;
      7'b0000001: n2402_o = n2401_o;
      default: n2402_o = n2400_o;
    endcase
  assign n2403_o = n2242_o[31:24];
  assign n2404_o = n2270_o[23:16];
  assign n2405_o = n2298_o[15:8];
  assign n2406_o = n2326_o[7:0];
  assign n2407_o = write_data_r[95:88];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2408_o = n2405_o;
      7'b0100000: n2408_o = n2404_o;
      7'b0010000: n2408_o = n2403_o;
      7'b0001000: n2408_o = n2407_o;
      7'b0000100: n2408_o = n2407_o;
      7'b0000010: n2408_o = n2407_o;
      7'b0000001: n2408_o = n2407_o;
      default: n2408_o = n2406_o;
    endcase
  assign n2409_o = n2270_o[31:24];
  assign n2410_o = n2298_o[23:16];
  assign n2411_o = n2326_o[15:8];
  assign n2412_o = write_data_r[103:96];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2413_o = n2410_o;
      7'b0100000: n2413_o = n2409_o;
      7'b0010000: n2413_o = n2412_o;
      7'b0001000: n2413_o = n2412_o;
      7'b0000100: n2413_o = n2412_o;
      7'b0000010: n2413_o = n2412_o;
      7'b0000001: n2413_o = n2412_o;
      default: n2413_o = n2411_o;
    endcase
  assign n2414_o = n2298_o[31:24];
  assign n2415_o = n2326_o[23:16];
  assign n2416_o = write_data_r[111:104];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2417_o = n2414_o;
      7'b0100000: n2417_o = n2416_o;
      7'b0010000: n2417_o = n2416_o;
      7'b0001000: n2417_o = n2416_o;
      7'b0000100: n2417_o = n2416_o;
      7'b0000010: n2417_o = n2416_o;
      7'b0000001: n2417_o = n2416_o;
      default: n2417_o = n2415_o;
    endcase
  assign n2418_o = n2326_o[31:24];
  assign n2419_o = write_data_r[119:112];
  /* ../../HW/src/top/ddr_tx.vhd:498:5  */
  always @*
    case (n2327_o)
      7'b1000000: n2420_o = n2419_o;
      7'b0100000: n2420_o = n2419_o;
      7'b0010000: n2420_o = n2419_o;
      7'b0001000: n2420_o = n2419_o;
      7'b0000100: n2420_o = n2419_o;
      7'b0000010: n2420_o = n2419_o;
      7'b0000001: n2420_o = n2419_o;
      default: n2420_o = n2418_o;
    endcase
  assign n2421_o = {n2420_o, n2417_o, n2413_o, n2408_o, n2402_o, n2395_o, n2387_o, n2378_o, n2369_o, n2360_o, n2352_o, n2345_o, n2339_o, n2334_o, n2330_o};
  assign n2422_o = write_data_r[119:0];
  /* ../../HW/src/top/ddr_tx.vhd:497:1  */
  assign n2423_o = write2 ? n2421_o : n2422_o;
  assign n2424_o = write_data_r[127:120];
  /* ../../HW/src/top/ddr_tx.vhd:585:13  */
  assign n2428_o = ~reset_in;
  /* ../../HW/src/top/ddr_tx.vhd:593:70  */
  assign n2430_o = byteenable[15:8];
  /* ../../HW/src/top/ddr_tx.vhd:595:65  */
  assign n2432_o = write_data[127:64];
  /* ../../HW/src/top/ddr_tx.vhd:596:38  */
  assign n2433_o = write_data[63:0];
  /* ../../HW/src/top/ddr_tx.vhd:598:8  */
  assign n2434_o = write2 ? write_data : write_data_r;
  /* ../../HW/src/top/ddr_tx.vhd:598:8  */
  assign n2435_o = write2 ? byteenable : byteenable_r;
  assign n2437_o = n2434_o[63:0];
  /* ../../HW/src/top/ddr_tx.vhd:592:8  */
  assign n2438_o = write_data_write_ena ? n2432_o : n2437_o;
  assign n2439_o = n2434_o[127:64];
  assign n2440_o = write_data_r[127:64];
  /* ../../HW/src/top/ddr_tx.vhd:592:8  */
  assign n2441_o = write_data_write_ena ? n2440_o : n2439_o;
  assign n2443_o = {8'b00000000, n2430_o};
  /* ../../HW/src/top/ddr_tx.vhd:592:8  */
  assign n2444_o = write_data_write_ena ? n2443_o : n2435_o;
  assign n2446_o = {n2441_o, n2438_o};
  /* ../../HW/src/top/ddr_tx.vhd:591:5  */
  assign n2459_o = write_data_write_ena ? write_data_write : write_data_write_r;
  /* ../../HW/src/top/ddr_tx.vhd:591:5  */
  always @(posedge clock_in or posedge n2428_o)
    if (n2428_o)
      n2460_q <= 41'b00000000000000000000000000000000000000000;
    else
      n2460_q <= n2459_o;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  assign n2461_o = n1707_o ? write_data_write_ena : write_data_write_ena_r;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  always @(posedge clock_in or posedge n1705_o)
    if (n1705_o)
      n2462_q <= 1'b0;
    else
      n2462_q <= n2461_o;
  assign n2466_o = {n2424_o, n2423_o};
  /* ../../HW/src/top/ddr_tx.vhd:591:5  */
  always @(posedge clock_in or posedge n2428_o)
    if (n2428_o)
      n2467_q <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n2467_q <= n2446_o;
  /* ../../HW/src/top/ddr_tx.vhd:591:5  */
  assign n2468_o = write_data_write_ena ? n2433_o : write_data_2_r;
  /* ../../HW/src/top/ddr_tx.vhd:591:5  */
  always @(posedge clock_in or posedge n2428_o)
    if (n2428_o)
      n2469_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n2469_q <= n2468_o;
  /* ../../HW/src/top/ddr_tx.vhd:591:5  */
  always @(posedge clock_in or posedge n2428_o)
    if (n2428_o)
      n2470_q <= 16'b0000000000000000;
    else
      n2470_q <= n2444_o;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  assign n2472_o = write_data_write_ena ? n1720_o : write_next_addr_r;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  always @(posedge clock_in or posedge n1705_o)
    if (n1705_o)
      n2473_q <= 32'b00000000000000000000000000000000;
    else
      n2473_q <= n2472_o;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  assign n2474_o = write_data_write_ena ? n1717_o : write_flush_r;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  always @(posedge clock_in or posedge n1705_o)
    if (n1705_o)
      n2475_q <= 1'b0;
    else
      n2475_q <= n2474_o;
  /* ../../HW/src/top/ddr_tx.vhd:230:9  */
  assign n2476_o = awvalid ? n1662_o : write_request_r;
  /* ../../HW/src/top/ddr_tx.vhd:230:9  */
  always @(posedge clock_in or posedge n1654_o)
    if (n1654_o)
      n2477_q <= 10'b0000000000;
    else
      n2477_q <= n2476_o;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  assign n2478_o = ddr_bresp_in ? n1723_o : write_complete_r;
  /* ../../HW/src/top/ddr_tx.vhd:283:7  */
  always @(posedge clock_in or posedge n1705_o)
    if (n1705_o)
      n2479_q <= 10'b0000000000;
    else
      n2479_q <= n2478_o;
  /* ../../HW/src/top/ddr_tx.vhd:230:9  */
  always @(posedge clock_in or posedge n1654_o)
    if (n1654_o)
      n2480_q <= 3'b000;
    else
      n2480_q <= n1668_o;
  /* ../../HW/src/top/ddr_tx.vhd:230:9  */
  assign n2481_o = n1658_o ? n1659_o : awaddr_r;
  /* ../../HW/src/top/ddr_tx.vhd:230:9  */
  always @(posedge clock_in or posedge n1654_o)
    if (n1654_o)
      n2482_q <= 32'b00000000000000000000000000000000;
    else
      n2482_q <= n2481_o;
endmodule

module ddr_rx
  (input  clock_in,
   input  reset_in,
   input  [31:0] read_addr_in,
   input  read_cs_in,
   input  read_in,
   input  read_vm_in,
   input  [2:0] read_vector_in,
   input  read_fork_in,
   input  [3:0] read_start_in,
   input  [3:0] read_end_in,
   input  read_data_wait_in,
   input  [4:0] read_burstlen_in,
   input  [15:0] read_filler_data_in,
   input  ddr_rvalid_in,
   input  ddr_rlast_in,
   input  [63:0] ddr_rdata_in,
   input  ddr_arready_in,
   output read_data_ready_out,
   output read_fork_out,
   output read_data_valid_out,
   output read_data_valid_vm_out,
   output [63:0] read_data_out,
   output read_wait_request_out,
   output [31:0] ddr_araddr_out,
   output [2:0] ddr_arlen_out,
   output ddr_arvalid_out,
   output ddr_rready_out,
   output [1:0] ddr_arburst_out,
   output [3:0] ddr_arcache_out,
   output ddr_arid_out,
   output ddr_arlock_out,
   output [2:0] ddr_arprot_out,
   output [3:0] ddr_arqos_out,
   output [2:0] ddr_arsize_out);
  wire [4:0] read_burstlen_r;
  wire [4:0] next_read_burstlen;
  wire burstbegin;
  wire read_data_valid;
  wire rvalid;
  wire [34:0] read_record_write;
  wire [34:0] read_record_write_r;
  wire read_record_write_ena;
  wire read_record_write_ena_r;
  wire read_record_read_ena;
  wire read_record_read_empty;
  wire read_record_read_full;
  wire read_record_read_full_r;
  wire [34:0] read_record_read;
  wire read_data_read_ena;
  wire read_data_read_ena_2;
  wire read_data_read_empty;
  wire [63:0] read_data_read;
  wire read_wait_request;
  wire [127:0] read_data_read_r;
  wire [1:0] read_data_read_valid_r;
  wire read_data_write_full;
  wire read2;
  wire ddr_read;
  wire [31:0] rd_ddr_addr;
  wire [4:0] rd_ddr_burstlen;
  wire read_data_ready;
  wire [4:0] read_burstlen2;
  wire [4:0] read_burstlen3;
  wire [31:0] read_addr;
  wire read_piggyback;
  wire read_piggyback_r;
  wire [63:0] read_data;
  wire read_pause_r;
  wire [31:0] read_pause_addr_r;
  wire [2:0] read_pause_burstlen_r;
  wire read_fifo_read_ena;
  wire read_fifo_read_empty;
  wire read_fifo_write_ena;
  wire read_fifo_write_full;
  wire [36:0] read_fifo_write;
  wire [36:0] read_fifo_read;
  wire [36:0] read_fifo_write_flat;
  wire [36:0] read_fifo_read_flat;
  wire [12:0] read_complete_r;
  wire [12:0] read_request_r;
  wire read_pending_full_r;
  wire [9:0] read_transaction_complete_r;
  wire [9:0] read_transaction_request_r;
  wire [63:0] read_data_fifo_i_n946;
  wire read_data_fifo_i_n949;
  wire read_data_fifo_i_n950;
  wire [63:0] read_data_fifo_i_q_out;
  wire [8:0] read_data_fifo_i_ravail_out;
  wire [8:0] read_data_fifo_i_wused_out;
  wire read_data_fifo_i_empty_out;
  wire read_data_fifo_i_full_out;
  wire read_data_fifo_i_almost_full_out;
  wire n962_o;
  wire n963_o;
  wire n964_o;
  wire n967_o;
  wire n968_o;
  wire n969_o;
  wire n972_o;
  wire n973_o;
  wire n974_o;
  wire n975_o;
  wire [36:0] ddr_rx_fifo_i_n977;
  wire ddr_rx_fifo_i_n980;
  wire ddr_rx_fifo_i_n981;
  wire [36:0] ddr_rx_fifo_i_q_out;
  wire [3:0] ddr_rx_fifo_i_ravail_out;
  wire [3:0] ddr_rx_fifo_i_wused_out;
  wire ddr_rx_fifo_i_empty_out;
  wire ddr_rx_fifo_i_full_out;
  wire ddr_rx_fifo_i_almost_full_out;
  wire [31:0] n999_o;
  wire [2:0] n1002_o;
  wire n1004_o;
  wire n1006_o;
  wire [36:0] n1007_o;
  wire [31:0] n1015_o;
  wire [2:0] n1018_o;
  wire [2:0] n1020_o;
  wire n1022_o;
  wire n1024_o;
  wire [36:0] n1025_o;
  wire [2:0] n1032_o;
  wire [31:0] n1033_o;
  wire [2:0] n1034_o;
  wire n1036_o;
  wire n1037_o;
  localparam n1042_o = 1'b0;
  localparam [1:0] n1043_o = 2'b01;
  localparam [3:0] n1044_o = 4'b0011;
  localparam n1045_o = 1'b0;
  localparam [2:0] n1046_o = 3'b000;
  localparam [3:0] n1047_o = 4'b0000;
  localparam [2:0] n1048_o = 3'b011;
  wire [31:0] n1051_o;
  wire [2:0] n1052_o;
  wire n1053_o;
  wire n1054_o;
  wire n1055_o;
  wire n1056_o;
  wire [34:0] read_record_fifo_i_n1058;
  wire read_record_fifo_i_n1061;
  wire read_record_fifo_i_n1063;
  wire [34:0] read_record_fifo_i_q_out;
  wire [5:0] read_record_fifo_i_ravail_out;
  wire [5:0] read_record_fifo_i_wused_out;
  wire read_record_fifo_i_empty_out;
  wire read_record_fifo_i_full_out;
  wire read_record_fifo_i_almost_full_out;
  wire n1073_o;
  wire n1074_o;
  wire n1075_o;
  wire n1076_o;
  wire n1077_o;
  wire n1078_o;
  wire n1079_o;
  wire n1080_o;
  wire n1081_o;
  wire n1082_o;
  wire n1083_o;
  wire n1084_o;
  wire n1086_o;
  wire n1087_o;
  wire n1088_o;
  wire n1089_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1095_o;
  wire n1096_o;
  wire n1098_o;
  wire n1099_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1108_o;
  wire n1109_o;
  wire [8:0] n1120_o;
  wire [2:0] n1121_o;
  wire [8:0] n1122_o;
  wire n1124_o;
  wire n1126_o;
  wire [8:0] n1128_o;
  wire [8:0] n1130_o;
  wire n1132_o;
  wire n1134_o;
  wire [8:0] n1136_o;
  wire [8:0] n1138_o;
  wire n1140_o;
  wire n1142_o;
  wire [8:0] n1144_o;
  wire [8:0] n1146_o;
  wire n1148_o;
  wire [8:0] n1150_o;
  wire [8:0] n1151_o;
  wire [8:0] n1152_o;
  wire [8:0] n1153_o;
  wire [8:0] n1154_o;
  wire [8:0] n1155_o;
  wire [8:0] n1156_o;
  wire [8:0] n1157_o;
  wire [8:0] n1159_o;
  wire [8:0] n1161_o;
  wire [4:0] n1162_o;
  wire [4:0] n1163_o;
  wire n1167_o;
  wire n1169_o;
  wire n1170_o;
  wire n1171_o;
  wire [2:0] n1172_o;
  wire n1173_o;
  wire n1175_o;
  wire n1177_o;
  wire [3:0] n1199_o;
  wire [3:0] n1200_o;
  wire [15:0] n1201_o;
  wire [3:0] n1203_o;
  wire n1205_o;
  wire n1207_o;
  wire n1208_o;
  wire [7:0] n1209_o;
  wire [7:0] n1210_o;
  wire [7:0] n1211_o;
  wire [3:0] n1213_o;
  wire n1215_o;
  wire n1217_o;
  wire n1218_o;
  wire [7:0] n1219_o;
  wire [7:0] n1220_o;
  wire [7:0] n1221_o;
  wire [3:0] n1223_o;
  wire n1225_o;
  wire n1227_o;
  wire n1228_o;
  wire [7:0] n1229_o;
  wire [7:0] n1230_o;
  wire [7:0] n1231_o;
  wire [3:0] n1233_o;
  wire n1235_o;
  wire n1237_o;
  wire n1238_o;
  wire [7:0] n1239_o;
  wire [7:0] n1240_o;
  wire [7:0] n1241_o;
  wire [3:0] n1243_o;
  wire n1245_o;
  wire n1247_o;
  wire n1248_o;
  wire [7:0] n1249_o;
  wire [7:0] n1250_o;
  wire [7:0] n1251_o;
  wire [3:0] n1253_o;
  wire n1255_o;
  wire n1257_o;
  wire n1258_o;
  wire [7:0] n1259_o;
  wire [7:0] n1260_o;
  wire [7:0] n1261_o;
  wire [3:0] n1263_o;
  wire n1265_o;
  wire n1267_o;
  wire n1268_o;
  wire [7:0] n1269_o;
  wire [7:0] n1270_o;
  wire [7:0] n1271_o;
  wire [3:0] n1273_o;
  wire n1275_o;
  wire n1277_o;
  wire n1278_o;
  wire [7:0] n1279_o;
  wire [7:0] n1280_o;
  wire [7:0] n1281_o;
  wire [2:0] n1286_o;
  wire [63:0] n1287_o;
  wire n1289_o;
  wire [63:0] n1290_o;
  wire n1292_o;
  wire [63:0] n1293_o;
  wire n1295_o;
  wire [63:0] n1296_o;
  wire n1298_o;
  wire [63:0] n1299_o;
  wire n1301_o;
  wire [63:0] n1302_o;
  wire n1304_o;
  wire [63:0] n1305_o;
  wire n1307_o;
  wire [63:0] n1308_o;
  wire [6:0] n1309_o;
  reg [63:0] n1310_o;
  wire [2:0] n1319_o;
  wire n1321_o;
  wire n1324_o;
  wire [2:0] n1325_o;
  wire [3:0] n1326_o;
  wire [3:0] n1327_o;
  wire [3:0] n1328_o;
  wire n1329_o;
  wire [2:0] n1330_o;
  wire [2:0] n1331_o;
  wire n1333_o;
  wire n1336_o;
  wire n1337_o;
  wire n1340_o;
  wire n1341_o;
  wire n1342_o;
  wire n1345_o;
  wire n1348_o;
  wire n1350_o;
  wire n1352_o;
  wire n1353_o;
  wire n1355_o;
  wire n1356_o;
  wire n1357_o;
  wire [28:0] n1364_o;
  wire n1366_o;
  wire [31:0] n1367_o;
  wire [4:0] n1369_o;
  wire [31:0] n1370_o;
  wire [31:0] n1372_o;
  wire [31:0] n1373_o;
  wire [4:0] n1374_o;
  wire n1380_o;
  wire n1381_o;
  wire [4:0] n1383_o;
  wire [4:0] n1384_o;
  wire n1385_o;
  wire [4:0] n1387_o;
  wire [4:0] n1388_o;
  wire [4:0] n1389_o;
  wire [4:0] n1390_o;
  wire n1394_o;
  wire n1419_o;
  wire n1420_o;
  wire n1421_o;
  wire n1422_o;
  wire n1423_o;
  wire n1424_o;
  wire n1425_o;
  wire n1426_o;
  wire n1430_o;
  wire [12:0] n1433_o;
  wire [2:0] n1435_o;
  wire [12:0] n1436_o;
  wire [12:0] n1437_o;
  wire [9:0] n1440_o;
  wire n1442_o;
  wire [9:0] n1444_o;
  wire [12:0] n1446_o;
  wire n1448_o;
  wire [9:0] n1449_o;
  wire n1451_o;
  wire n1452_o;
  wire n1455_o;
  wire n1456_o;
  wire n1457_o;
  wire n1458_o;
  wire n1460_o;
  wire [63:0] n1461_o;
  wire n1462_o;
  wire n1463_o;
  wire [127:0] n1464_o;
  wire [63:0] n1465_o;
  wire [63:0] n1466_o;
  wire [63:0] n1467_o;
  wire [63:0] n1468_o;
  wire [63:0] n1469_o;
  wire [1:0] n1470_o;
  wire [1:0] n1471_o;
  wire [1:0] n1472_o;
  wire n1473_o;
  wire n1474_o;
  wire [63:0] n1475_o;
  wire n1476_o;
  wire n1477_o;
  wire n1478_o;
  wire n1479_o;
  wire n1480_o;
  wire [63:0] n1481_o;
  wire [63:0] n1482_o;
  wire n1483_o;
  wire n1484_o;
  wire [127:0] n1485_o;
  wire [63:0] n1486_o;
  wire [63:0] n1487_o;
  wire [63:0] n1488_o;
  wire [63:0] n1489_o;
  wire [63:0] n1490_o;
  wire [1:0] n1491_o;
  wire n1492_o;
  wire n1493_o;
  wire n1494_o;
  wire n1495_o;
  wire n1496_o;
  wire [127:0] n1497_o;
  wire [127:0] n1498_o;
  wire [127:0] n1499_o;
  wire [1:0] n1500_o;
  wire [1:0] n1501_o;
  reg [4:0] n1525_q;
  wire [34:0] n1526_o;
  reg [34:0] n1527_q;
  reg n1528_q;
  reg n1532_q;
  reg [127:0] n1533_q;
  reg [1:0] n1534_q;
  wire n1536_o;
  reg n1537_q;
  reg n1538_q;
  wire [31:0] n1539_o;
  reg [31:0] n1540_q;
  wire [2:0] n1541_o;
  reg [2:0] n1542_q;
  wire [36:0] n1543_o;
  wire [12:0] n1544_o;
  reg [12:0] n1545_q;
  wire [12:0] n1546_o;
  reg [12:0] n1547_q;
  reg n1548_q;
  wire [9:0] n1549_o;
  reg [9:0] n1550_q;
  wire [9:0] n1551_o;
  reg [9:0] n1552_q;
  wire [63:0] n1553_o;
  assign read_data_ready_out = read_data_ready;
  assign read_fork_out = n1074_o;
  assign read_data_valid_out = read_data_valid;
  assign read_data_valid_vm_out = n1073_o;
  assign read_data_out = n1553_o;
  assign read_wait_request_out = read_wait_request;
  assign ddr_araddr_out = n1051_o;
  assign ddr_arlen_out = n1052_o;
  assign ddr_arvalid_out = n1055_o;
  assign ddr_rready_out = n1056_o;
  assign ddr_arburst_out = n1043_o;
  assign ddr_arcache_out = n1044_o;
  assign ddr_arid_out = n1042_o;
  assign ddr_arlock_out = n1045_o;
  assign ddr_arprot_out = n1046_o;
  assign ddr_arqos_out = n1047_o;
  assign ddr_arsize_out = n1048_o;
  /* ../../HW/src/top/ddr_rx.vhd:156:8  */
  assign read_burstlen_r = n1525_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:157:8  */
  assign next_read_burstlen = n1390_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:158:8  */
  assign burstbegin = n1105_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:159:8  */
  assign read_data_valid = n1084_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:160:8  */
  assign rvalid = n964_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:162:8  */
  assign read_record_write = n1526_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:163:8  */
  assign read_record_write_r = n1527_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:164:8  */
  assign read_record_write_ena = n1357_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:165:8  */
  assign read_record_write_ena_r = n1528_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:168:8  */
  assign read_record_read_ena = read_data_valid; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:169:8  */
  assign read_record_read_empty = read_record_fifo_i_n1061; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:171:8  */
  assign read_record_read_full = read_record_fifo_i_n1063; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:172:8  */
  assign read_record_read_full_r = n1532_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:173:8  */
  assign read_record_read = read_record_fifo_i_n1058; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:175:8  */
  assign read_data_read_ena = n1092_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:176:8  */
  assign read_data_read_ena_2 = n1426_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:177:8  */
  assign read_data_read_empty = read_data_fifo_i_n949; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:178:8  */
  assign read_data_read = read_data_fifo_i_n946; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:179:8  */
  assign read_wait_request = n1096_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:181:8  */
  assign read_data_read_r = n1533_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:182:8  */
  assign read_data_read_valid_r = n1534_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:183:8  */
  assign read_data_write_full = read_data_fifo_i_n950; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:185:8  */
  assign read2 = n1099_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:187:8  */
  assign ddr_read = n1109_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:190:8  */
  assign rd_ddr_addr = n1373_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:191:8  */
  assign rd_ddr_burstlen = n1374_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:192:8  */
  assign read_data_ready = n1082_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:194:8  */
  assign read_burstlen2 = n1163_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:195:8  */
  assign read_burstlen3 = n1162_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:196:8  */
  assign read_addr = read_addr_in; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:198:8  */
  assign read_piggyback = n1355_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:199:8  */
  assign read_piggyback_r = n1537_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:201:8  */
  assign read_data = n1310_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:202:8  */
  assign read_pause_r = n1538_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:203:8  */
  assign read_pause_addr_r = n1540_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:204:8  */
  assign read_pause_burstlen_r = n1542_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:206:8  */
  assign read_fifo_read_ena = n969_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:207:8  */
  assign read_fifo_read_empty = ddr_rx_fifo_i_n980; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:208:8  */
  assign read_fifo_write_ena = n975_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:209:8  */
  assign read_fifo_write_full = ddr_rx_fifo_i_n981; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:210:8  */
  assign read_fifo_write = n1543_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:211:8  */
  assign read_fifo_read = n1007_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:212:8  */
  assign read_fifo_write_flat = n1025_o; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:213:8  */
  assign read_fifo_read_flat = ddr_rx_fifo_i_n977; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:218:8  */
  assign read_complete_r = n1545_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:219:8  */
  assign read_request_r = n1547_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:220:8  */
  assign read_pending_full_r = n1548_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:222:8  */
  assign read_transaction_complete_r = n1550_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:223:8  */
  assign read_transaction_request_r = n1552_q; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:247:16  */
  assign read_data_fifo_i_n946 = read_data_fifo_i_q_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:250:20  */
  assign read_data_fifo_i_n949 = read_data_fifo_i_empty_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:251:19  */
  assign read_data_fifo_i_n950 = read_data_fifo_i_full_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:233:1  */
  scfifo_64_9_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 read_data_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(ddr_rdata_in),
    .write_in(rvalid),
    .read_in(read_data_read_ena_2),
    .q_out(read_data_fifo_i_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(read_data_fifo_i_empty_out),
    .full_out(read_data_fifo_i_full_out),
    .almost_full_out());
  /* ../../HW/src/top/ddr_rx.vhd:256:63  */
  assign n962_o = ~read_data_write_full;
  /* ../../HW/src/top/ddr_rx.vhd:256:39  */
  assign n963_o = n962_o & ddr_rvalid_in;
  /* ../../HW/src/top/ddr_rx.vhd:256:15  */
  assign n964_o = n963_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:258:54  */
  assign n967_o = ~read_fifo_read_empty;
  /* ../../HW/src/top/ddr_rx.vhd:258:60  */
  assign n968_o = ddr_arready_in & n967_o;
  /* ../../HW/src/top/ddr_rx.vhd:258:27  */
  assign n969_o = n968_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:260:49  */
  assign n972_o = read_fifo_write[35];
  /* ../../HW/src/top/ddr_rx.vhd:260:82  */
  assign n973_o = ~read_fifo_write_full;
  /* ../../HW/src/top/ddr_rx.vhd:260:58  */
  assign n974_o = n973_o & n972_o;
  /* ../../HW/src/top/ddr_rx.vhd:260:28  */
  assign n975_o = n974_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:281:16  */
  assign ddr_rx_fifo_i_n977 = ddr_rx_fifo_i_q_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:284:20  */
  assign ddr_rx_fifo_i_n980 = ddr_rx_fifo_i_empty_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:285:19  */
  assign ddr_rx_fifo_i_n981 = ddr_rx_fifo_i_full_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:267:1  */
  scfifo_37_4_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 ddr_rx_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(read_fifo_write_flat),
    .write_in(read_fifo_write_ena),
    .read_in(read_fifo_read_ena),
    .q_out(ddr_rx_fifo_i_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(ddr_rx_fifo_i_empty_out),
    .full_out(ddr_rx_fifo_i_full_out),
    .almost_full_out());
  /* ../../HW/src/top/ddr_rx.vhd:132:22  */
  assign n999_o = read_fifo_read_flat[36:5];
  /* ../../HW/src/top/ddr_rx.vhd:134:35  */
  assign n1002_o = read_fifo_read_flat[4:2];
  /* ../../HW/src/top/ddr_rx.vhd:136:22  */
  assign n1004_o = read_fifo_read_flat[1];
  /* ../../HW/src/top/ddr_rx.vhd:138:28  */
  assign n1006_o = read_fifo_read_flat[0];
  /* ../../HW/src/top/ztachip.vhd:595:1  */
  assign n1007_o = {n1006_o, n1004_o, n1002_o, n999_o};
  /* ../../HW/src/top/ddr_rx.vhd:112:81  */
  assign n1015_o = read_fifo_write[31:0];
  /* ../../HW/src/top/ddr_rx.vhd:114:102  */
  assign n1018_o = read_fifo_write[34:32];
  /* ../../HW/src/top/ddr_rx.vhd:114:110  */
  assign n1020_o = n1018_o - 3'b001;
  /* ../../HW/src/top/ddr_rx.vhd:116:38  */
  assign n1022_o = read_fifo_write[35];
  /* ../../HW/src/top/ddr_rx.vhd:118:38  */
  assign n1024_o = read_fifo_write[36];
  /* ../../HW/src/top/ztachip.vhd:676:30  */
  assign n1025_o = {n1015_o, n1020_o, n1022_o, n1024_o};
  /* ../../HW/src/top/ddr_rx.vhd:308:36  */
  assign n1032_o = rd_ddr_burstlen[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:302:4  */
  assign n1033_o = read_pause_r ? read_pause_addr_r : rd_ddr_addr;
  /* ../../HW/src/top/ddr_rx.vhd:302:4  */
  assign n1034_o = read_pause_r ? read_pause_burstlen_r : n1032_o;
  /* ../../HW/src/top/ddr_rx.vhd:302:4  */
  assign n1036_o = read_pause_r ? 1'b1 : ddr_read;
  /* ../../HW/src/top/ddr_rx.vhd:311:32  */
  assign n1037_o = burstbegin & ddr_read;
  /* ../../HW/src/top/ddr_rx.vhd:335:37  */
  assign n1051_o = read_fifo_read[31:0];
  /* ../../HW/src/top/ddr_rx.vhd:336:36  */
  assign n1052_o = read_fifo_read[34:32];
  /* ../../HW/src/top/ddr_rx.vhd:337:38  */
  assign n1053_o = read_fifo_read[36];
  /* ../../HW/src/top/ddr_rx.vhd:337:54  */
  assign n1054_o = ~read_fifo_read_empty;
  /* ../../HW/src/top/ddr_rx.vhd:337:49  */
  assign n1055_o = n1053_o & n1054_o;
  /* ../../HW/src/top/ddr_rx.vhd:338:23  */
  assign n1056_o = ~read_data_write_full;
  /* ../../HW/src/top/ddr_rx.vhd:360:16  */
  assign read_record_fifo_i_n1058 = read_record_fifo_i_q_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:363:20  */
  assign read_record_fifo_i_n1061 = read_record_fifo_i_empty_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:365:26  */
  assign read_record_fifo_i_n1063 = read_record_fifo_i_almost_full_out; // (signal)
  /* ../../HW/src/top/ddr_rx.vhd:345:1  */
  scfifo_35_6_53_bf8b4530d8d246dd74ac53a13471bba17941dff7 read_record_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(read_record_write_r),
    .write_in(read_record_write_ena_r),
    .read_in(read_record_read_ena),
    .q_out(read_record_fifo_i_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(read_record_fifo_i_empty_out),
    .full_out(),
    .almost_full_out(read_record_fifo_i_almost_full_out));
  /* ../../HW/src/top/ddr_rx.vhd:374:43  */
  assign n1073_o = read_record_read[18];
  /* ../../HW/src/top/ddr_rx.vhd:375:34  */
  assign n1074_o = read_record_read[17];
  /* ../../HW/src/top/ddr_rx.vhd:376:43  */
  assign n1075_o = read_data_read_valid_r[1];
  /* ../../HW/src/top/ddr_rx.vhd:376:74  */
  assign n1076_o = read_data_read_valid_r[0];
  /* ../../HW/src/top/ddr_rx.vhd:376:102  */
  assign n1077_o = read_record_read[7];
  /* ../../HW/src/top/ddr_rx.vhd:376:82  */
  assign n1078_o = ~n1077_o;
  /* ../../HW/src/top/ddr_rx.vhd:376:78  */
  assign n1079_o = n1076_o | n1078_o;
  /* ../../HW/src/top/ddr_rx.vhd:376:47  */
  assign n1080_o = n1075_o & n1079_o;
  /* ../../HW/src/top/ddr_rx.vhd:376:154  */
  assign n1081_o = ~read_record_read_empty;
  /* ../../HW/src/top/ddr_rx.vhd:376:149  */
  assign n1082_o = n1080_o & n1081_o;
  /* ../../HW/src/top/ddr_rx.vhd:377:41  */
  assign n1083_o = ~read_data_wait_in;
  /* ../../HW/src/top/ddr_rx.vhd:377:36  */
  assign n1084_o = read_data_ready & n1083_o;
  /* ../../HW/src/top/ddr_rx.vhd:383:35  */
  assign n1086_o = read_record_read[3];
  /* ../../HW/src/top/ddr_rx.vhd:384:35  */
  assign n1087_o = read_record_read[7];
  /* ../../HW/src/top/ddr_rx.vhd:383:60  */
  assign n1088_o = n1086_o | n1087_o;
  /* ../../HW/src/top/ddr_rx.vhd:385:35  */
  assign n1089_o = read_record_read[8];
  /* ../../HW/src/top/ddr_rx.vhd:384:81  */
  assign n1090_o = n1088_o | n1089_o;
  /* ../../HW/src/top/ddr_rx.vhd:381:39  */
  assign n1091_o = n1090_o & read_data_valid;
  /* ../../HW/src/top/ddr_rx.vhd:380:27  */
  assign n1092_o = n1091_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:391:61  */
  assign n1095_o = read_record_read_full_r | read_pause_r;
  /* ../../HW/src/top/ddr_rx.vhd:391:26  */
  assign n1096_o = n1095_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:393:41  */
  assign n1098_o = ~read_wait_request;
  /* ../../HW/src/top/ddr_rx.vhd:393:18  */
  assign n1099_o = n1098_o ? read_in : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:399:54  */
  assign n1103_o = read_burstlen_r == 5'b00000;
  /* ../../HW/src/top/ddr_rx.vhd:399:35  */
  assign n1104_o = n1103_o & read2;
  /* ../../HW/src/top/ddr_rx.vhd:399:19  */
  assign n1105_o = n1104_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:401:38  */
  assign n1108_o = read2 & burstbegin;
  /* ../../HW/src/top/ddr_rx.vhd:401:17  */
  assign n1109_o = n1108_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:417:18  */
  assign n1120_o = {4'b0, read_burstlen_in};  //  uext
  /* ../../HW/src/top/ddr_rx.vhd:418:39  */
  assign n1121_o = read_addr[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:418:14  */
  assign n1122_o = {6'b0, n1121_o};  //  uext
  /* ../../HW/src/top/ddr_rx.vhd:419:31  */
  assign n1124_o = read_vector_in == 3'b001;
  /* ../../HW/src/top/ddr_rx.vhd:420:21  */
  assign n1126_o = $unsigned(n1120_o) > $unsigned(9'b000010100);
  /* ../../HW/src/top/ddr_rx.vhd:420:7  */
  assign n1128_o = n1126_o ? 9'b000010100 : n1120_o;
  /* ../../HW/src/top/ddr_rx.vhd:423:28  */
  assign n1130_o = n1128_o << 32'b00000000000000000000000000000001;
  /* ../../HW/src/top/ddr_rx.vhd:424:34  */
  assign n1132_o = read_vector_in == 3'b011;
  /* ../../HW/src/top/ddr_rx.vhd:425:21  */
  assign n1134_o = $unsigned(n1120_o) > $unsigned(9'b000001010);
  /* ../../HW/src/top/ddr_rx.vhd:425:7  */
  assign n1136_o = n1134_o ? 9'b000001010 : n1120_o;
  /* ../../HW/src/top/ddr_rx.vhd:428:28  */
  assign n1138_o = n1136_o << 32'b00000000000000000000000000000010;
  /* ../../HW/src/top/ddr_rx.vhd:429:34  */
  assign n1140_o = read_vector_in == 3'b111;
  /* ../../HW/src/top/ddr_rx.vhd:430:21  */
  assign n1142_o = $unsigned(n1120_o) > $unsigned(9'b000000101);
  /* ../../HW/src/top/ddr_rx.vhd:430:7  */
  assign n1144_o = n1142_o ? 9'b000000101 : n1120_o;
  /* ../../HW/src/top/ddr_rx.vhd:433:28  */
  assign n1146_o = n1144_o << 32'b00000000000000000000000000000011;
  /* ../../HW/src/top/ddr_rx.vhd:435:21  */
  assign n1148_o = $unsigned(n1120_o) > $unsigned(9'b000101000);
  /* ../../HW/src/top/ddr_rx.vhd:435:7  */
  assign n1150_o = n1148_o ? 9'b000101000 : n1120_o;
  /* ../../HW/src/top/ddr_rx.vhd:429:4  */
  assign n1151_o = n1140_o ? n1144_o : n1150_o;
  /* ../../HW/src/top/ddr_rx.vhd:429:4  */
  assign n1152_o = n1140_o ? n1146_o : n1150_o;
  /* ../../HW/src/top/ddr_rx.vhd:424:4  */
  assign n1153_o = n1132_o ? n1136_o : n1151_o;
  /* ../../HW/src/top/ddr_rx.vhd:424:4  */
  assign n1154_o = n1132_o ? n1138_o : n1152_o;
  /* ../../HW/src/top/ddr_rx.vhd:419:4  */
  assign n1155_o = n1124_o ? n1128_o : n1153_o;
  /* ../../HW/src/top/ddr_rx.vhd:419:4  */
  assign n1156_o = n1124_o ? n1130_o : n1154_o;
  /* ../../HW/src/top/ddr_rx.vhd:440:21  */
  assign n1157_o = n1156_o + n1122_o;
  /* ../../HW/src/top/ddr_rx.vhd:440:28  */
  assign n1159_o = n1157_o + 9'b000000111;
  /* ../../HW/src/top/ddr_rx.vhd:441:23  */
  assign n1161_o = n1159_o >> 32'b00000000000000000000000000000011;
  /* ../../HW/src/top/ddr_rx.vhd:442:22  */
  assign n1162_o = n1161_o[4:0];  // trunc
  /* ../../HW/src/top/ddr_rx.vhd:443:22  */
  assign n1163_o = n1155_o[4:0];  // trunc
  /* ../../HW/src/top/ddr_rx.vhd:448:17  */
  assign n1167_o = ~reset_in;
  /* ../../HW/src/top/ddr_rx.vhd:455:61  */
  assign n1169_o = read_record_read_full | read_pending_full_r;
  /* ../../HW/src/top/ddr_rx.vhd:456:30  */
  assign n1170_o = read_fifo_write_full & burstbegin;
  /* ../../HW/src/top/ddr_rx.vhd:456:59  */
  assign n1171_o = ddr_read & n1170_o;
  /* ../../HW/src/top/ddr_rx.vhd:458:55  */
  assign n1172_o = rd_ddr_burstlen[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:460:38  */
  assign n1173_o = ~read_fifo_write_full;
  /* ../../HW/src/top/ddr_rx.vhd:460:12  */
  assign n1175_o = n1173_o ? 1'b0 : read_pause_r;
  /* ../../HW/src/top/ddr_rx.vhd:456:12  */
  assign n1177_o = n1171_o ? 1'b1 : n1175_o;
  /* ../../HW/src/top/ddr_rx.vhd:483:38  */
  assign n1199_o = read_record_read[12:9];
  /* ../../HW/src/top/ddr_rx.vhd:484:38  */
  assign n1200_o = read_record_read[16:13];
  /* ../../HW/src/top/ddr_rx.vhd:486:32  */
  assign n1201_o = read_record_read[34:19];
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1203_o = n1199_o + 4'b0000;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1205_o = $signed(n1203_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1207_o = $unsigned(n1200_o) > $unsigned(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1208_o = n1207_o & n1205_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1209_o = read_data[7:0];
  /* ../../HW/src/top/ddr_rx.vhd:493:82  */
  assign n1210_o = n1201_o[7:0];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1211_o = n1208_o ? n1209_o : n1210_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1213_o = n1199_o + 4'b0001;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1215_o = $signed(n1213_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1217_o = $unsigned(n1200_o) > $unsigned(4'b0001);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1218_o = n1217_o & n1215_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1219_o = read_data[15:8];
  /* ../../HW/src/top/ddr_rx.vhd:495:82  */
  assign n1220_o = n1201_o[15:8];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1221_o = n1218_o ? n1219_o : n1220_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1223_o = n1199_o + 4'b0010;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1225_o = $signed(n1223_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1227_o = $unsigned(n1200_o) > $unsigned(4'b0010);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1228_o = n1227_o & n1225_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1229_o = read_data[23:16];
  /* ../../HW/src/top/ddr_rx.vhd:493:82  */
  assign n1230_o = n1201_o[7:0];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1231_o = n1228_o ? n1229_o : n1230_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1233_o = n1199_o + 4'b0011;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1235_o = $signed(n1233_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1237_o = $unsigned(n1200_o) > $unsigned(4'b0011);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1238_o = n1237_o & n1235_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1239_o = read_data[31:24];
  /* ../../HW/src/top/ddr_rx.vhd:495:82  */
  assign n1240_o = n1201_o[15:8];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1241_o = n1238_o ? n1239_o : n1240_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1243_o = n1199_o + 4'b0100;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1245_o = $signed(n1243_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1247_o = $unsigned(n1200_o) > $unsigned(4'b0100);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1248_o = n1247_o & n1245_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1249_o = read_data[39:32];
  /* ../../HW/src/top/ddr_rx.vhd:493:82  */
  assign n1250_o = n1201_o[7:0];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1251_o = n1248_o ? n1249_o : n1250_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1253_o = n1199_o + 4'b0101;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1255_o = $signed(n1253_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1257_o = $unsigned(n1200_o) > $unsigned(4'b0101);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1258_o = n1257_o & n1255_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1259_o = read_data[47:40];
  /* ../../HW/src/top/ddr_rx.vhd:495:82  */
  assign n1260_o = n1201_o[15:8];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1261_o = n1258_o ? n1259_o : n1260_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1263_o = n1199_o + 4'b0110;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1265_o = $signed(n1263_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1267_o = $unsigned(n1200_o) > $unsigned(4'b0110);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1268_o = n1267_o & n1265_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1269_o = read_data[55:48];
  /* ../../HW/src/top/ddr_rx.vhd:493:82  */
  assign n1270_o = n1201_o[7:0];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1271_o = n1268_o ? n1269_o : n1270_o;
  /* ../../HW/src/top/ddr_rx.vhd:488:17  */
  assign n1273_o = n1199_o + 4'b0111;
  /* ../../HW/src/top/ddr_rx.vhd:488:52  */
  assign n1275_o = $signed(n1273_o) >= $signed(4'b0000);
  /* ../../HW/src/top/ddr_rx.vhd:489:16  */
  assign n1277_o = $unsigned(n1200_o) > $unsigned(4'b0111);
  /* ../../HW/src/top/ddr_rx.vhd:488:57  */
  assign n1278_o = n1277_o & n1275_o;
  /* ../../HW/src/top/ddr_rx.vhd:490:80  */
  assign n1279_o = read_data[63:56];
  /* ../../HW/src/top/ddr_rx.vhd:495:82  */
  assign n1280_o = n1201_o[15:8];
  /* ../../HW/src/top/ddr_rx.vhd:488:7  */
  assign n1281_o = n1278_o ? n1279_o : n1280_o;
  /* ../../HW/src/top/ddr_rx.vhd:507:26  */
  assign n1286_o = read_record_read[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:509:71  */
  assign n1287_o = read_data_read_r[63:0];
  /* ../../HW/src/top/ddr_rx.vhd:508:9  */
  assign n1289_o = n1286_o == 3'b000;
  /* ../../HW/src/top/ddr_rx.vhd:511:71  */
  assign n1290_o = read_data_read_r[71:8];
  /* ../../HW/src/top/ddr_rx.vhd:510:9  */
  assign n1292_o = n1286_o == 3'b001;
  /* ../../HW/src/top/ddr_rx.vhd:513:71  */
  assign n1293_o = read_data_read_r[79:16];
  /* ../../HW/src/top/ddr_rx.vhd:512:9  */
  assign n1295_o = n1286_o == 3'b010;
  /* ../../HW/src/top/ddr_rx.vhd:515:71  */
  assign n1296_o = read_data_read_r[87:24];
  /* ../../HW/src/top/ddr_rx.vhd:514:9  */
  assign n1298_o = n1286_o == 3'b011;
  /* ../../HW/src/top/ddr_rx.vhd:517:71  */
  assign n1299_o = read_data_read_r[95:32];
  /* ../../HW/src/top/ddr_rx.vhd:516:9  */
  assign n1301_o = n1286_o == 3'b100;
  /* ../../HW/src/top/ddr_rx.vhd:519:71  */
  assign n1302_o = read_data_read_r[103:40];
  /* ../../HW/src/top/ddr_rx.vhd:518:9  */
  assign n1304_o = n1286_o == 3'b101;
  /* ../../HW/src/top/ddr_rx.vhd:521:71  */
  assign n1305_o = read_data_read_r[111:48];
  /* ../../HW/src/top/ddr_rx.vhd:520:9  */
  assign n1307_o = n1286_o == 3'b110;
  /* ../../HW/src/top/ddr_rx.vhd:523:71  */
  assign n1308_o = read_data_read_r[119:56];
  assign n1309_o = {n1307_o, n1304_o, n1301_o, n1298_o, n1295_o, n1292_o, n1289_o};
  /* ../../HW/src/top/ddr_rx.vhd:507:5  */
  always @*
    case (n1309_o)
      7'b1000000: n1310_o = n1305_o;
      7'b0100000: n1310_o = n1302_o;
      7'b0010000: n1310_o = n1299_o;
      7'b0001000: n1310_o = n1296_o;
      7'b0000100: n1310_o = n1293_o;
      7'b0000010: n1310_o = n1290_o;
      7'b0000001: n1310_o = n1287_o;
      default: n1310_o = n1308_o;
    endcase
  /* ../../HW/src/top/ddr_rx.vhd:535:65  */
  assign n1319_o = read_addr[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:536:25  */
  assign n1321_o = next_read_burstlen == 5'b00000;
  /* ../../HW/src/top/ddr_rx.vhd:536:4  */
  assign n1324_o = n1321_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:541:37  */
  assign n1325_o = read_addr[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:541:12  */
  assign n1326_o = {1'b0, n1325_o};  //  uext
  /* ../../HW/src/top/ddr_rx.vhd:542:12  */
  assign n1327_o = {1'b0, read_vector_in};  //  uext
  /* ../../HW/src/top/ddr_rx.vhd:541:91  */
  assign n1328_o = n1326_o + n1327_o;
  /* ../../HW/src/top/ddr_rx.vhd:544:22  */
  assign n1329_o = n1328_o[3];
  /* ../../HW/src/top/ddr_rx.vhd:546:26  */
  assign n1330_o = read_addr[2:0];
  /* ../../HW/src/top/ddr_rx.vhd:546:58  */
  assign n1331_o = n1330_o + read_vector_in;
  /* ../../HW/src/top/ddr_rx.vhd:546:83  */
  assign n1333_o = n1331_o == 3'b111;
  /* ../../HW/src/top/ddr_rx.vhd:546:4  */
  assign n1336_o = n1333_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:552:21  */
  assign n1337_o = ~n1324_o;
  /* ../../HW/src/top/ddr_rx.vhd:556:27  */
  assign n1340_o = $unsigned(read_burstlen_in) > $unsigned(5'b00001);
  /* ../../HW/src/top/ddr_rx.vhd:559:42  */
  assign n1341_o = ~n1336_o;
  /* ../../HW/src/top/ddr_rx.vhd:559:26  */
  assign n1342_o = n1329_o | n1341_o;
  /* ../../HW/src/top/ddr_rx.vhd:559:10  */
  assign n1345_o = n1342_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/ddr_rx.vhd:559:10  */
  assign n1348_o = n1342_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:556:7  */
  assign n1350_o = n1340_o ? n1345_o : 1'b1;
  /* ../../HW/src/top/ddr_rx.vhd:556:7  */
  assign n1352_o = n1340_o ? n1348_o : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:552:4  */
  assign n1353_o = n1337_o ? 1'b0 : n1350_o;
  /* ../../HW/src/top/ddr_rx.vhd:552:4  */
  assign n1355_o = n1337_o ? 1'b0 : n1352_o;
  /* ../../HW/src/top/ddr_rx.vhd:586:40  */
  assign n1356_o = ~read_wait_request;
  /* ../../HW/src/top/ddr_rx.vhd:586:35  */
  assign n1357_o = read2 & n1356_o;
  /* ../../HW/src/top/ddr_rx.vhd:599:125  */
  assign n1364_o = read_addr[31:3];
  /* ../../HW/src/top/ddr_rx.vhd:601:23  */
  assign n1366_o = ~read_piggyback_r;
  assign n1367_o = {n1364_o, 3'b000};
  /* ../../HW/src/top/ddr_rx.vhd:605:50  */
  assign n1369_o = read_burstlen3 - 5'b00001;
  assign n1370_o = {n1364_o, 3'b000};
  /* ../../HW/src/top/ddr_rx.vhd:606:60  */
  assign n1372_o = n1370_o + 32'b00000000000000000000000000001000;
  /* ../../HW/src/top/ddr_rx.vhd:601:4  */
  assign n1373_o = n1366_o ? n1367_o : n1372_o;
  /* ../../HW/src/top/ddr_rx.vhd:601:4  */
  assign n1374_o = n1366_o ? read_burstlen3 : n1369_o;
  /* ../../HW/src/top/ddr_rx.vhd:619:22  */
  assign n1380_o = read_burstlen_r == 5'b00000;
  /* ../../HW/src/top/ddr_rx.vhd:620:27  */
  assign n1381_o = ~read_wait_request;
  /* ../../HW/src/top/ddr_rx.vhd:621:46  */
  assign n1383_o = read_burstlen2 - 5'b00001;
  /* ../../HW/src/top/ddr_rx.vhd:620:7  */
  assign n1384_o = n1381_o ? n1383_o : read_burstlen_r;
  /* ../../HW/src/top/ddr_rx.vhd:626:27  */
  assign n1385_o = ~read_wait_request;
  /* ../../HW/src/top/ddr_rx.vhd:627:47  */
  assign n1387_o = read_burstlen_r - 5'b00001;
  /* ../../HW/src/top/ddr_rx.vhd:626:7  */
  assign n1388_o = n1385_o ? n1387_o : read_burstlen_r;
  /* ../../HW/src/top/ddr_rx.vhd:619:4  */
  assign n1389_o = n1380_o ? n1384_o : n1388_o;
  /* ../../HW/src/top/ddr_rx.vhd:618:1  */
  assign n1390_o = read2 ? n1389_o : read_burstlen_r;
  /* ../../HW/src/top/ddr_rx.vhd:640:17  */
  assign n1394_o = ~reset_in;
  /* ../../HW/src/top/ddr_rx.vhd:664:26  */
  assign n1419_o = ~read_data_read_empty;
  /* ../../HW/src/top/ddr_rx.vhd:664:105  */
  assign n1420_o = read_data_read_valid_r[1];
  /* ../../HW/src/top/ddr_rx.vhd:664:108  */
  assign n1421_o = ~n1420_o;
  /* ../../HW/src/top/ddr_rx.vhd:664:80  */
  assign n1422_o = read_data_read_ena | n1421_o;
  /* ../../HW/src/top/ddr_rx.vhd:664:138  */
  assign n1423_o = read_data_read_valid_r[0];
  /* ../../HW/src/top/ddr_rx.vhd:664:141  */
  assign n1424_o = ~n1423_o;
  /* ../../HW/src/top/ddr_rx.vhd:664:113  */
  assign n1425_o = n1422_o | n1424_o;
  /* ../../HW/src/top/ddr_rx.vhd:664:52  */
  assign n1426_o = n1425_o ? n1419_o : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:668:13  */
  assign n1430_o = ~reset_in;
  /* ../../HW/src/top/ddr_rx.vhd:682:45  */
  assign n1433_o = read_complete_r + 13'b0000000000001;
  /* ../../HW/src/top/ddr_rx.vhd:685:67  */
  assign n1435_o = read_fifo_write[34:32];
  /* ../../HW/src/top/ddr_rx.vhd:685:44  */
  assign n1436_o = {10'b0, n1435_o};  //  uext
  /* ../../HW/src/top/ddr_rx.vhd:685:43  */
  assign n1437_o = read_request_r + n1436_o;
  /* ../../HW/src/top/ddr_rx.vhd:689:67  */
  assign n1440_o = read_transaction_request_r + 10'b0000000001;
  /* ../../HW/src/top/ddr_rx.vhd:691:22  */
  assign n1442_o = ddr_rlast_in & rvalid;
  /* ../../HW/src/top/ddr_rx.vhd:692:69  */
  assign n1444_o = read_transaction_complete_r + 10'b0000000001;
  /* ../../HW/src/top/ddr_rx.vhd:694:35  */
  assign n1446_o = read_request_r - read_complete_r;
  /* ../../HW/src/top/ddr_rx.vhd:694:61  */
  assign n1448_o = $signed(n1446_o) >= $signed(13'b0000111110110);
  /* ../../HW/src/top/ddr_rx.vhd:695:47  */
  assign n1449_o = read_transaction_request_r - read_transaction_complete_r;
  /* ../../HW/src/top/ddr_rx.vhd:695:85  */
  assign n1451_o = $signed(n1449_o) >= $signed(10'b0000111111);
  /* ../../HW/src/top/ddr_rx.vhd:694:140  */
  assign n1452_o = n1448_o | n1451_o;
  /* ../../HW/src/top/ddr_rx.vhd:694:8  */
  assign n1455_o = n1452_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ddr_rx.vhd:702:30  */
  assign n1456_o = read_record_read[3];
  /* ../../HW/src/top/ddr_rx.vhd:702:75  */
  assign n1457_o = read_record_read[7];
  /* ../../HW/src/top/ddr_rx.vhd:702:55  */
  assign n1458_o = n1457_o & n1456_o;
  /* ../../HW/src/top/ddr_rx.vhd:705:43  */
  assign n1460_o = ~read_data_read_empty;
  /* ../../HW/src/top/ddr_rx.vhd:709:79  */
  assign n1461_o = read_data_read_r[127:64];
  /* ../../HW/src/top/ddr_rx.vhd:710:65  */
  assign n1462_o = read_data_read_valid_r[0];
  /* ../../HW/src/top/ddr_rx.vhd:712:43  */
  assign n1463_o = ~read_data_read_empty;
  assign n1464_o = {read_data_read, n1461_o};
  assign n1465_o = n1464_o[63:0];
  assign n1466_o = read_data_read_r[63:0];
  /* ../../HW/src/top/ddr_rx.vhd:702:11  */
  assign n1467_o = n1458_o ? n1466_o : n1465_o;
  assign n1468_o = n1464_o[127:64];
  /* ../../HW/src/top/ddr_rx.vhd:702:11  */
  assign n1469_o = n1458_o ? read_data_read : n1468_o;
  assign n1470_o = {n1462_o, n1463_o};
  assign n1471_o = {1'b0, n1460_o};
  /* ../../HW/src/top/ddr_rx.vhd:702:11  */
  assign n1472_o = n1458_o ? n1471_o : n1470_o;
  /* ../../HW/src/top/ddr_rx.vhd:715:36  */
  assign n1473_o = read_data_read_valid_r[1];
  /* ../../HW/src/top/ddr_rx.vhd:715:39  */
  assign n1474_o = ~n1473_o;
  /* ../../HW/src/top/ddr_rx.vhd:716:79  */
  assign n1475_o = read_data_read_r[127:64];
  /* ../../HW/src/top/ddr_rx.vhd:717:65  */
  assign n1476_o = read_data_read_valid_r[0];
  /* ../../HW/src/top/ddr_rx.vhd:718:43  */
  assign n1477_o = ~read_data_read_empty;
  /* ../../HW/src/top/ddr_rx.vhd:720:39  */
  assign n1478_o = read_data_read_valid_r[0];
  /* ../../HW/src/top/ddr_rx.vhd:720:42  */
  assign n1479_o = ~n1478_o;
  /* ../../HW/src/top/ddr_rx.vhd:721:43  */
  assign n1480_o = ~read_data_read_empty;
  assign n1481_o = read_data_read_r[127:64];
  /* ../../HW/src/top/ddr_rx.vhd:720:11  */
  assign n1482_o = n1479_o ? read_data_read : n1481_o;
  assign n1483_o = read_data_read_valid_r[0];
  /* ../../HW/src/top/ddr_rx.vhd:720:11  */
  assign n1484_o = n1479_o ? n1480_o : n1483_o;
  assign n1485_o = {read_data_read, n1475_o};
  assign n1486_o = n1485_o[63:0];
  assign n1487_o = read_data_read_r[63:0];
  /* ../../HW/src/top/ddr_rx.vhd:715:11  */
  assign n1488_o = n1474_o ? n1486_o : n1487_o;
  assign n1489_o = n1485_o[127:64];
  /* ../../HW/src/top/ddr_rx.vhd:715:11  */
  assign n1490_o = n1474_o ? n1489_o : n1482_o;
  assign n1491_o = {n1476_o, n1477_o};
  assign n1492_o = n1491_o[0];
  /* ../../HW/src/top/ddr_rx.vhd:715:11  */
  assign n1493_o = n1474_o ? n1492_o : n1484_o;
  assign n1494_o = n1491_o[1];
  assign n1495_o = read_data_read_valid_r[1];
  /* ../../HW/src/top/ddr_rx.vhd:715:11  */
  assign n1496_o = n1474_o ? n1494_o : n1495_o;
  assign n1497_o = {n1490_o, n1488_o};
  assign n1498_o = {n1469_o, n1467_o};
  /* ../../HW/src/top/ddr_rx.vhd:701:8  */
  assign n1499_o = read_data_read_ena ? n1498_o : n1497_o;
  assign n1500_o = {n1496_o, n1493_o};
  /* ../../HW/src/top/ddr_rx.vhd:701:8  */
  assign n1501_o = read_data_read_ena ? n1472_o : n1500_o;
  /* ../../HW/src/top/ddr_rx.vhd:649:9  */
  always @(posedge clock_in or posedge n1394_o)
    if (n1394_o)
      n1525_q <= 5'b00000;
    else
      n1525_q <= next_read_burstlen;
  /* ../../HW/src/top/ddr_rx.vhd:640:5  */
  assign n1526_o = {read_filler_data_in, read_vm_in, read_fork_in, read_end_in, read_start_in, n1336_o, n1329_o, read_vector_in, n1353_o, n1319_o};
  /* ../../HW/src/top/ddr_rx.vhd:649:9  */
  always @(posedge clock_in or posedge n1394_o)
    if (n1394_o)
      n1527_q <= 35'b00000000000000000000000000000000000;
    else
      n1527_q <= read_record_write;
  /* ../../HW/src/top/ddr_rx.vhd:649:9  */
  always @(posedge clock_in or posedge n1394_o)
    if (n1394_o)
      n1528_q <= 1'b0;
    else
      n1528_q <= read_record_write_ena;
  /* ../../HW/src/top/ddr_rx.vhd:454:9  */
  always @(posedge clock_in or posedge n1167_o)
    if (n1167_o)
      n1532_q <= 1'b0;
    else
      n1532_q <= n1169_o;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1533_q <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n1533_q <= n1499_o;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1534_q <= 2'b00;
    else
      n1534_q <= n1501_o;
  /* ../../HW/src/top/ddr_rx.vhd:649:9  */
  assign n1536_o = read_record_write_ena ? read_piggyback : read_piggyback_r;
  /* ../../HW/src/top/ddr_rx.vhd:649:9  */
  always @(posedge clock_in or posedge n1394_o)
    if (n1394_o)
      n1537_q <= 1'b0;
    else
      n1537_q <= n1536_o;
  /* ../../HW/src/top/ddr_rx.vhd:454:9  */
  always @(posedge clock_in or posedge n1167_o)
    if (n1167_o)
      n1538_q <= 1'b0;
    else
      n1538_q <= n1177_o;
  /* ../../HW/src/top/ddr_rx.vhd:454:9  */
  assign n1539_o = n1171_o ? rd_ddr_addr : read_pause_addr_r;
  /* ../../HW/src/top/ddr_rx.vhd:454:9  */
  always @(posedge clock_in or posedge n1167_o)
    if (n1167_o)
      n1540_q <= 32'b00000000000000000000000000000000;
    else
      n1540_q <= n1539_o;
  /* ../../HW/src/top/ddr_rx.vhd:454:9  */
  assign n1541_o = n1171_o ? n1172_o : read_pause_burstlen_r;
  /* ../../HW/src/top/ddr_rx.vhd:454:9  */
  always @(posedge clock_in or posedge n1167_o)
    if (n1167_o)
      n1542_q <= 3'b000;
    else
      n1542_q <= n1541_o;
  /* ../../HW/src/top/ddr_rx.vhd:448:5  */
  assign n1543_o = {n1037_o, n1036_o, n1034_o, n1033_o};
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  assign n1544_o = read_data_read_ena_2 ? n1433_o : read_complete_r;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1545_q <= 13'b0000000000000;
    else
      n1545_q <= n1544_o;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  assign n1546_o = read_fifo_write_ena ? n1437_o : read_request_r;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1547_q <= 13'b0000000000000;
    else
      n1547_q <= n1546_o;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1548_q <= 1'b0;
    else
      n1548_q <= n1455_o;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  assign n1549_o = n1442_o ? n1444_o : read_transaction_complete_r;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1550_q <= 10'b0000000000;
    else
      n1550_q <= n1549_o;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  assign n1551_o = read_fifo_write_ena ? n1440_o : read_transaction_request_r;
  /* ../../HW/src/top/ddr_rx.vhd:677:5  */
  always @(posedge clock_in or posedge n1430_o)
    if (n1430_o)
      n1552_q <= 10'b0000000000;
    else
      n1552_q <= n1551_o;
  /* ../../HW/src/top/ddr_rx.vhd:668:1  */
  assign n1553_o = {n1281_o, n1271_o, n1261_o, n1251_o, n1241_o, n1231_o, n1221_o, n1211_o};
endmodule

module sram_core
  (input  clock_in,
   input  reset_in,
   input  [14:0] dp_rd_addr_in,
   input  [14:0] dp_wr_addr_in,
   input  dp_rd_fork_in,
   input  dp_wr_fork_in,
   input  dp_write_in,
   input  [2:0] dp_write_vector_in,
   input  dp_read_in,
   input  dp_read_vm_in,
   input  [2:0] dp_read_vector_in,
   input  dp_read_gen_valid_in,
   input  [63:0] dp_writedata_in,
   output dp_readdatavalid_out,
   output dp_readdatavalid_vm_out,
   output [63:0] dp_readdata_out);
  wire [1:0] write;
  wire [1:0] read;
  wire [63:0] writedata;
  wire [1:0] readdatavalid;
  wire [127:0] readdata;
  wire vm_r;
  wire vm_rr;
  wire vm_rrr;
  wire vm_rrrr;
  wire n852_o;
  wire n853_o;
  wire n857_o;
  wire n860_o;
  reg n862_o;
  reg n863_o;
  reg [63:0] n864_o;
  wire n868_o;
  wire n871_o;
  reg n873_o;
  reg n874_o;
  wire n878_o;
  wire [63:0] n879_o;
  wire [63:0] n880_o;
  wire [63:0] n881_o;
  wire n885_o;
  wire [13:0] n900_o;
  wire [13:0] n901_o;
  wire n902_o;
  wire n903_o;
  wire gen_sram_n1_sram_i_n904;
  wire [63:0] gen_sram_n1_sram_i_n905;
  wire gen_sram_n1_sram_i_dp_readdatavalid_out;
  wire [63:0] gen_sram_n1_sram_i_dp_readdata_out;
  wire [13:0] n910_o;
  wire [13:0] n911_o;
  wire n912_o;
  wire n913_o;
  wire gen_sram_n2_sram_i_n914;
  wire [63:0] gen_sram_n2_sram_i_n915;
  wire gen_sram_n2_sram_i_dp_readdatavalid_out;
  wire [63:0] gen_sram_n2_sram_i_dp_readdata_out;
  wire [1:0] n920_o;
  wire [1:0] n921_o;
  wire [1:0] n922_o;
  wire [127:0] n923_o;
  reg n924_q;
  reg n925_q;
  reg n926_q;
  reg n927_q;
  assign dp_readdatavalid_out = n853_o;
  assign dp_readdatavalid_vm_out = vm_rrrr;
  assign dp_readdata_out = n881_o;
  /* ../../HW/src/top/sram_core.vhd:55:8  */
  assign write = n920_o; // (signal)
  /* ../../HW/src/top/sram_core.vhd:56:8  */
  assign read = n921_o; // (signal)
  /* ../../HW/src/top/sram_core.vhd:57:8  */
  assign writedata = n864_o; // (signal)
  /* ../../HW/src/top/sram_core.vhd:58:8  */
  assign readdatavalid = n922_o; // (signal)
  /* ../../HW/src/top/sram_core.vhd:59:8  */
  assign readdata = n923_o; // (signal)
  /* ../../HW/src/top/sram_core.vhd:60:8  */
  assign vm_r = n924_q; // (signal)
  /* ../../HW/src/top/sram_core.vhd:61:8  */
  assign vm_rr = n925_q; // (signal)
  /* ../../HW/src/top/sram_core.vhd:62:8  */
  assign vm_rrr = n926_q; // (signal)
  /* ../../HW/src/top/sram_core.vhd:63:8  */
  assign vm_rrrr = n927_q; // (signal)
  /* ../../HW/src/top/sram_core.vhd:66:47  */
  assign n852_o = readdatavalid == 2'b00;
  /* ../../HW/src/top/sram_core.vhd:66:29  */
  assign n853_o = n852_o ? 1'b0 : 1'b1;
  /* ../../HW/src/top/sram_core.vhd:73:22  */
  assign n857_o = dp_wr_addr_in[14];
  /* ../../HW/src/top/sram_core.vhd:74:7  */
  assign n860_o = n857_o == 1'b0;
  /* ../../HW/src/top/sram_core.vhd:73:4  */
  always @*
    case (n860_o)
      1'b1: n862_o = dp_write_in;
      default: n862_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram_core.vhd:73:4  */
  always @*
    case (n860_o)
      1'b1: n863_o = 1'b0;
      default: n863_o = dp_write_in;
    endcase
  /* ../../HW/src/top/sram_core.vhd:73:4  */
  always @*
    case (n860_o)
      1'b1: n864_o = dp_writedata_in;
      default: n864_o = dp_writedata_in;
    endcase
  /* ../../HW/src/top/sram_core.vhd:89:22  */
  assign n868_o = dp_rd_addr_in[14];
  /* ../../HW/src/top/sram_core.vhd:90:7  */
  assign n871_o = n868_o == 1'b0;
  /* ../../HW/src/top/sram_core.vhd:89:4  */
  always @*
    case (n871_o)
      1'b1: n873_o = dp_read_in;
      default: n873_o = 1'b0;
    endcase
  /* ../../HW/src/top/sram_core.vhd:89:4  */
  always @*
    case (n871_o)
      1'b1: n874_o = 1'b0;
      default: n874_o = dp_read_in;
    endcase
  /* ../../HW/src/top/sram_core.vhd:103:17  */
  assign n878_o = readdatavalid[0];
  /* ../../HW/src/top/sram_core.vhd:104:60  */
  assign n879_o = readdata[63:0];
  /* ../../HW/src/top/sram_core.vhd:106:60  */
  assign n880_o = readdata[127:64];
  /* ../../HW/src/top/sram_core.vhd:103:1  */
  assign n881_o = n878_o ? n879_o : n880_o;
  /* ../../HW/src/top/sram_core.vhd:113:17  */
  assign n885_o = ~reset_in;
  /* ../../HW/src/top/sram_core.vhd:137:39  */
  assign n900_o = dp_rd_addr_in[13:0];
  /* ../../HW/src/top/sram_core.vhd:138:39  */
  assign n901_o = dp_wr_addr_in[13:0];
  /* ../../HW/src/top/sram_core.vhd:139:29  */
  assign n902_o = write[0];
  /* ../../HW/src/top/sram_core.vhd:141:25  */
  assign n903_o = read[0];
  /* ../../HW/src/top/sram_core.vhd:145:31  */
  assign gen_sram_n1_sram_i_n904 = gen_sram_n1_sram_i_dp_readdatavalid_out; // (signal)
  /* ../../HW/src/top/sram_core.vhd:146:28  */
  assign gen_sram_n1_sram_i_n905 = gen_sram_n1_sram_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/sram_core.vhd:130:1  */
  sram_14 gen_sram_n1_sram_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .dp_rd_addr_in(n900_o),
    .dp_wr_addr_in(n901_o),
    .dp_write_in(n902_o),
    .dp_write_vector_in(dp_write_vector_in),
    .dp_read_in(n903_o),
    .dp_read_vector_in(dp_read_vector_in),
    .dp_read_gen_valid_in(dp_read_gen_valid_in),
    .dp_writedata_in(writedata),
    .dp_readdatavalid_out(gen_sram_n1_sram_i_dp_readdatavalid_out),
    .dp_readdata_out(gen_sram_n1_sram_i_dp_readdata_out));
  /* ../../HW/src/top/sram_core.vhd:137:39  */
  assign n910_o = dp_rd_addr_in[13:0];
  /* ../../HW/src/top/sram_core.vhd:138:39  */
  assign n911_o = dp_wr_addr_in[13:0];
  /* ../../HW/src/top/sram_core.vhd:139:29  */
  assign n912_o = write[1];
  /* ../../HW/src/top/sram_core.vhd:141:25  */
  assign n913_o = read[1];
  /* ../../HW/src/top/sram_core.vhd:145:31  */
  assign gen_sram_n2_sram_i_n914 = gen_sram_n2_sram_i_dp_readdatavalid_out; // (signal)
  /* ../../HW/src/top/sram_core.vhd:146:28  */
  assign gen_sram_n2_sram_i_n915 = gen_sram_n2_sram_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/sram_core.vhd:130:1  */
  sram_14 gen_sram_n2_sram_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .dp_rd_addr_in(n910_o),
    .dp_wr_addr_in(n911_o),
    .dp_write_in(n912_o),
    .dp_write_vector_in(dp_write_vector_in),
    .dp_read_in(n913_o),
    .dp_read_vector_in(dp_read_vector_in),
    .dp_read_gen_valid_in(dp_read_gen_valid_in),
    .dp_writedata_in(writedata),
    .dp_readdatavalid_out(gen_sram_n2_sram_i_dp_readdatavalid_out),
    .dp_readdata_out(gen_sram_n2_sram_i_dp_readdata_out));
  /* ../../HW/src/top/ztachip.vhd:540:23  */
  assign n920_o = {n863_o, n862_o};
  /* ../../HW/src/top/ztachip.vhd:539:26  */
  assign n921_o = {n874_o, n873_o};
  /* ../../HW/src/top/ztachip.vhd:538:26  */
  assign n922_o = {gen_sram_n2_sram_i_n914, gen_sram_n1_sram_i_n904};
  /* ../../HW/src/top/ztachip.vhd:537:25  */
  assign n923_o = {gen_sram_n2_sram_i_n915, gen_sram_n1_sram_i_n905};
  /* ../../HW/src/top/sram_core.vhd:119:9  */
  always @(posedge clock_in or posedge n885_o)
    if (n885_o)
      n924_q <= 1'b0;
    else
      n924_q <= dp_read_vm_in;
  /* ../../HW/src/top/sram_core.vhd:119:9  */
  always @(posedge clock_in or posedge n885_o)
    if (n885_o)
      n925_q <= 1'b0;
    else
      n925_q <= vm_r;
  /* ../../HW/src/top/sram_core.vhd:119:9  */
  always @(posedge clock_in or posedge n885_o)
    if (n885_o)
      n926_q <= 1'b0;
    else
      n926_q <= vm_rr;
  /* ../../HW/src/top/sram_core.vhd:119:9  */
  always @(posedge clock_in or posedge n885_o)
    if (n885_o)
      n927_q <= 1'b0;
    else
      n927_q <= vm_rrr;
endmodule

module axilite
  (input  clock_in,
   input  reset_in,
   input  [23:0] axilite_araddr_in,
   input  axilite_arvalid_in,
   input  axilite_rready_in,
   input  [23:0] axilite_awaddr_in,
   input  axilite_awvalid_in,
   input  axilite_wvalid_in,
   input  [31:0] axilite_wdata_in,
   input  axilite_bready_in,
   input  [31:0] bus_readdata_in,
   input  bus_readdatavalid_in,
   input  bus_writewait_in,
   input  bus_readwait_in,
   output axilite_arready_out,
   output axilite_rvalid_out,
   output axilite_rlast_out,
   output [31:0] axilite_rdata_out,
   output [1:0] axilite_rresp_out,
   output axilite_awready_out,
   output axilite_wready_out,
   output axilite_bvalid_out,
   output [1:0] axilite_bresp_out,
   output [23:0] bus_waddr_out,
   output [23:0] bus_raddr_out,
   output bus_write_out,
   output bus_read_out,
   output [31:0] bus_writedata_out);
  wire [31:0] axilite_rdata;
  wire bus_read;
  wire bus_readdatavalid_r;
  wire [31:0] bus_readdata_r;
  wire waddr_fifo_write;
  wire waddr_fifo_read;
  wire wdata_fifo_write;
  wire wdata_fifo_read;
  wire wdata_fifo_empty;
  wire wdata_fifo_full;
  wire waddr_fifo_empty;
  wire waddr_fifo_full;
  wire bus_write;
  wire n772_o;
  wire n773_o;
  wire [31:0] n774_o;
  wire n775_o;
  wire n777_o;
  wire n778_o;
  wire n779_o;
  wire n780_o;
  wire n781_o;
  wire n783_o;
  wire n784_o;
  localparam [1:0] n785_o = 2'b00;
  localparam [1:0] n786_o = 2'b00;
  wire n787_o;
  wire n788_o;
  wire n789_o;
  wire n790_o;
  wire [23:0] waddr_fifo_i_n791;
  wire waddr_fifo_i_n794;
  wire waddr_fifo_i_n795;
  wire [23:0] waddr_fifo_i_q_out;
  wire [5:0] waddr_fifo_i_ravail_out;
  wire [5:0] waddr_fifo_i_wused_out;
  wire waddr_fifo_i_empty_out;
  wire waddr_fifo_i_full_out;
  wire waddr_fifo_i_almost_full_out;
  wire n806_o;
  wire n807_o;
  wire n808_o;
  wire n809_o;
  wire [31:0] wdata_fifo_i_n810;
  wire wdata_fifo_i_n813;
  wire wdata_fifo_i_n814;
  wire [31:0] wdata_fifo_i_q_out;
  wire [5:0] wdata_fifo_i_ravail_out;
  wire [5:0] wdata_fifo_i_wused_out;
  wire wdata_fifo_i_empty_out;
  wire wdata_fifo_i_full_out;
  wire wdata_fifo_i_almost_full_out;
  wire n827_o;
  wire n829_o;
  wire n830_o;
  wire n831_o;
  wire n833_o;
  wire n835_o;
  reg n844_q;
  wire [31:0] n845_o;
  reg [31:0] n846_q;
  assign axilite_arready_out = n775_o;
  assign axilite_rvalid_out = n773_o;
  assign axilite_rlast_out = n772_o;
  assign axilite_rdata_out = axilite_rdata;
  assign axilite_rresp_out = n785_o;
  assign axilite_awready_out = n783_o;
  assign axilite_wready_out = n784_o;
  assign axilite_bvalid_out = waddr_fifo_read;
  assign axilite_bresp_out = n786_o;
  assign bus_waddr_out = waddr_fifo_i_n791;
  assign bus_raddr_out = axilite_araddr_in;
  assign bus_write_out = bus_write;
  assign bus_read_out = bus_read;
  assign bus_writedata_out = wdata_fifo_i_n810;
  /* ../../HW/src/top/axilite.vhd:66:8  */
  assign axilite_rdata = n774_o; // (signal)
  /* ../../HW/src/top/axilite.vhd:67:8  */
  assign bus_read = axilite_arvalid_in; // (signal)
  /* ../../HW/src/top/axilite.vhd:68:8  */
  assign bus_readdatavalid_r = n844_q; // (signal)
  /* ../../HW/src/top/axilite.vhd:69:8  */
  assign bus_readdata_r = n846_q; // (signal)
  /* ../../HW/src/top/axilite.vhd:70:8  */
  assign waddr_fifo_write = n788_o; // (signal)
  /* ../../HW/src/top/axilite.vhd:71:8  */
  assign waddr_fifo_read = n790_o; // (signal)
  /* ../../HW/src/top/axilite.vhd:72:8  */
  assign wdata_fifo_write = n807_o; // (signal)
  /* ../../HW/src/top/axilite.vhd:73:8  */
  assign wdata_fifo_read = n809_o; // (signal)
  /* ../../HW/src/top/axilite.vhd:74:8  */
  assign wdata_fifo_empty = wdata_fifo_i_n813; // (signal)
  /* ../../HW/src/top/axilite.vhd:75:8  */
  assign wdata_fifo_full = wdata_fifo_i_n814; // (signal)
  /* ../../HW/src/top/axilite.vhd:76:8  */
  assign waddr_fifo_empty = waddr_fifo_i_n794; // (signal)
  /* ../../HW/src/top/axilite.vhd:77:8  */
  assign waddr_fifo_full = waddr_fifo_i_n795; // (signal)
  /* ../../HW/src/top/axilite.vhd:78:8  */
  assign bus_write = n781_o; // (signal)
  /* ../../HW/src/top/axilite.vhd:87:43  */
  assign n772_o = bus_readdatavalid_in | bus_readdatavalid_r;
  /* ../../HW/src/top/axilite.vhd:89:44  */
  assign n773_o = bus_readdatavalid_in | bus_readdatavalid_r;
  /* ../../HW/src/top/axilite.vhd:91:34  */
  assign n774_o = bus_readdatavalid_in ? bus_readdata_in : bus_readdata_r;
  /* ../../HW/src/top/axilite.vhd:93:25  */
  assign n775_o = ~bus_readwait_in;
  /* ../../HW/src/top/axilite.vhd:97:40  */
  assign n777_o = ~waddr_fifo_empty;
  /* ../../HW/src/top/axilite.vhd:97:67  */
  assign n778_o = ~wdata_fifo_empty;
  /* ../../HW/src/top/axilite.vhd:97:46  */
  assign n779_o = n778_o & n777_o;
  /* ../../HW/src/top/axilite.vhd:97:73  */
  assign n780_o = axilite_bready_in & n779_o;
  /* ../../HW/src/top/axilite.vhd:97:18  */
  assign n781_o = n780_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/axilite.vhd:102:24  */
  assign n783_o = ~waddr_fifo_full;
  /* ../../HW/src/top/axilite.vhd:104:23  */
  assign n784_o = ~wdata_fifo_full;
  /* ../../HW/src/top/axilite.vhd:114:45  */
  assign n787_o = ~waddr_fifo_full;
  /* ../../HW/src/top/axilite.vhd:114:40  */
  assign n788_o = axilite_awvalid_in & n787_o;
  /* ../../HW/src/top/axilite.vhd:116:21  */
  assign n789_o = ~bus_writewait_in;
  /* ../../HW/src/top/axilite.vhd:116:43  */
  assign n790_o = n789_o & bus_write;
  /* ../../HW/src/top/axilite.vhd:132:16  */
  assign waddr_fifo_i_n791 = waddr_fifo_i_q_out; // (signal)
  /* ../../HW/src/top/axilite.vhd:135:20  */
  assign waddr_fifo_i_n794 = waddr_fifo_i_empty_out; // (signal)
  /* ../../HW/src/top/axilite.vhd:136:19  */
  assign waddr_fifo_i_n795 = waddr_fifo_i_full_out; // (signal)
  /* ../../HW/src/top/axilite.vhd:118:1  */
  scfifo_24_6_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 waddr_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(axilite_awaddr_in),
    .write_in(waddr_fifo_write),
    .read_in(waddr_fifo_read),
    .q_out(waddr_fifo_i_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(waddr_fifo_i_empty_out),
    .full_out(waddr_fifo_i_full_out),
    .almost_full_out());
  /* ../../HW/src/top/axilite.vhd:142:44  */
  assign n806_o = ~wdata_fifo_full;
  /* ../../HW/src/top/axilite.vhd:142:39  */
  assign n807_o = axilite_wvalid_in & n806_o;
  /* ../../HW/src/top/axilite.vhd:144:21  */
  assign n808_o = ~bus_writewait_in;
  /* ../../HW/src/top/axilite.vhd:144:43  */
  assign n809_o = n808_o & bus_write;
  /* ../../HW/src/top/axilite.vhd:160:16  */
  assign wdata_fifo_i_n810 = wdata_fifo_i_q_out; // (signal)
  /* ../../HW/src/top/axilite.vhd:163:20  */
  assign wdata_fifo_i_n813 = wdata_fifo_i_empty_out; // (signal)
  /* ../../HW/src/top/axilite.vhd:164:19  */
  assign wdata_fifo_i_n814 = wdata_fifo_i_full_out; // (signal)
  /* ../../HW/src/top/axilite.vhd:146:1  */
  scfifo_32_6_1_bf8b4530d8d246dd74ac53a13471bba17941dff7 wdata_fifo_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .data_in(axilite_wdata_in),
    .write_in(wdata_fifo_write),
    .read_in(wdata_fifo_read),
    .q_out(wdata_fifo_i_q_out),
    .ravail_out(),
    .wused_out(),
    .empty_out(wdata_fifo_i_empty_out),
    .full_out(wdata_fifo_i_full_out),
    .almost_full_out());
  /* ../../HW/src/top/axilite.vhd:172:16  */
  assign n827_o = ~reset_in;
  /* ../../HW/src/top/axilite.vhd:177:59  */
  assign n829_o = ~axilite_rready_in;
  /* ../../HW/src/top/axilite.vhd:177:38  */
  assign n830_o = n829_o & bus_readdatavalid_in;
  /* ../../HW/src/top/axilite.vhd:180:40  */
  assign n831_o = axilite_rready_in & bus_readdatavalid_r;
  /* ../../HW/src/top/axilite.vhd:180:10  */
  assign n833_o = n831_o ? 1'b0 : bus_readdatavalid_r;
  /* ../../HW/src/top/axilite.vhd:177:10  */
  assign n835_o = n830_o ? 1'b1 : n833_o;
  /* ../../HW/src/top/axilite.vhd:176:7  */
  always @(posedge clock_in or posedge n827_o)
    if (n827_o)
      n844_q <= 1'b0;
    else
      n844_q <= n835_o;
  /* ../../HW/src/top/axilite.vhd:176:7  */
  assign n845_o = n830_o ? bus_readdata_in : bus_readdata_r;
  /* ../../HW/src/top/axilite.vhd:176:7  */
  always @(posedge clock_in or posedge n827_o)
    if (n827_o)
      n846_q <= 32'b00000000000000000000000000000000;
    else
      n846_q <= n845_o;
endmodule

module ztachip
  (input  clock_in,
   input  clock_x2_in,
   input  reset_in,
   input  axi_rvalid_in,
   input  axi_rlast_in,
   input  [63:0] axi_rdata_in,
   input  axi_arready_in,
   input  axi_awready_in,
   input  axi_wready_in,
   input  axi_bresp_in,
   input  [23:0] axilite_araddr_in,
   input  axilite_arvalid_in,
   input  axilite_rready_in,
   input  [23:0] axilite_awaddr_in,
   input  axilite_awvalid_in,
   input  axilite_wvalid_in,
   input  [31:0] axilite_wdata_in,
   input  axilite_bready_in,
   output [31:0] axi_araddr_out,
   output [2:0] axi_arlen_out,
   output axi_arvalid_out,
   output axi_rready_out,
   output [1:0] axi_arburst_out,
   output [3:0] axi_arcache_out,
   output axi_arid_out,
   output axi_arlock_out,
   output [2:0] axi_arprot_out,
   output [3:0] axi_arqos_out,
   output [2:0] axi_arsize_out,
   output [31:0] axi_awaddr_out,
   output [2:0] axi_awlen_out,
   output axi_awvalid_out,
   output [31:0] axi_waddr_out,
   output axi_wvalid_out,
   output [63:0] axi_wdata_out,
   output axi_wlast_out,
   output [7:0] axi_wbe_out,
   output [1:0] axi_awburst_out,
   output [3:0] axi_awcache_out,
   output axi_awid_out,
   output axi_awlock_out,
   output [2:0] axi_awprot_out,
   output [3:0] axi_awqos_out,
   output [2:0] axi_awsize_out,
   output axi_bready_out,
   output axilite_arready_out,
   output axilite_rvalid_out,
   output axilite_rlast_out,
   output [31:0] axilite_rdata_out,
   output [1:0] axilite_rresp_out,
   output axilite_awready_out,
   output axilite_wready_out,
   output axilite_bvalid_out,
   output [1:0] axilite_bresp_out);
  wire [23:0] host_waddr;
  wire [23:0] host_raddr;
  wire host_wren;
  wire host_rden;
  wire [31:0] host_writedata;
  wire [31:0] host_readdata;
  wire host_readdatavalid;
  wire host_writewait;
  wire host_readwait;
  wire [1:0] pcore_busy;
  wire [1:0] busy;
  wire pcore_read_busy;
  wire pcore_write_busy;
  wire ready;
  wire [21:0] pcore_read_addr;
  wire pcore_read_fork;
  wire pcore_read_addr_mode;
  wire pcore_read_enable;
  wire pcore_read_gen_valid;
  wire [63:0] pcore_read_data;
  wire pcore_readdata_vm;
  wire pcore_read_data_valid;
  wire pcore_read_data_valid2;
  wire pcore_read_gen_valid2;
  wire [21:0] pcore_write_addr;
  wire pcore_write_fork;
  wire pcore_write_addr_mode;
  wire [5:0] pcore_mcast;
  wire pcore_write_enable;
  wire pcore_write_gen_valid;
  wire [63:0] pcore_write_data;
  wire [14:0] sram_read_addr;
  wire sram_read_fork;
  wire sram_read_enable;
  wire [2:0] sram_read_vector;
  wire sram_read_gen_valid;
  wire [63:0] sram_read_data;
  wire sram_read_data_valid;
  wire sram_readdata_vm;
  wire sram_read_vm;
  wire [14:0] sram_write_addr;
  wire sram_write_fork;
  wire sram_write_enable;
  wire [2:0] sram_write_vector;
  wire [63:0] sram_write_data;
  wire [31:0] ddr_read_addr;
  wire ddr_read_enable;
  wire ddr_read_enable_2;
  wire ddr_read_wait;
  wire ddr_read_wait_2;
  wire [63:0] ddr_read_data;
  wire ddr_read_data_valid;
  wire [4:0] ddr_read_burstlen;
  wire [15:0] ddr_read_filler_data;
  wire [31:0] ddr_write_addr;
  wire ddr_write_enable;
  wire ddr_write_enable_2;
  wire ddr_write_wait;
  wire ddr_write_wait_2;
  wire [63:0] ddr_write_data;
  wire [4:0] ddr_write_burstlen;
  wire [8:0] ddr_write_burstlen2;
  wire [4:0] ddr_write_burstlen3;
  wire ddr_data_ready;
  wire ddr_data_wait;
  wire [3:0] ddr_write_end;
  wire ddr_read_vm;
  wire ddr_readdata_vm;
  wire [10:0] task_start_addr;
  wire \task ;
  wire task_vm;
  wire [4:0] task_pcore;
  wire [71:0] bar;
  wire [47:0] pcore_write_counter_r;
  wire [47:0] sram_write_counter_r;
  wire [23:0] ddr_write_counter_r;
  wire dp_sram_read_fork;
  wire dp_sram_read_wait;
  wire dp_sram_write_fork;
  wire dp_sram_write_wait;
  wire dp_sram_write_enable;
  wire [2:0] dp_sram_write_vector;
  wire [17:0] dp_sram_write_addr;
  wire [63:0] dp_sram_write_data;
  wire [1:0] dp_sram_write_page;
  wire dp_sram_write_vm;
  wire dp_pcore_read_wait;
  wire dp_pcore_write_wait;
  wire [21:0] dp_pcore_write_addr;
  wire dp_pcore_write_fork;
  wire [63:0] dp_pcore_write_data;
  wire dp_pcore_write_enable;
  wire dp_pcore_write_vm;
  wire dp_pcore_read_vm;
  wire [21:0] dp_pcore_read_addr;
  wire dp_pcore_read_fork;
  wire dp_pcore_read_addr_mode;
  wire [17:0] dp_sram_read_addr;
  wire dp_pcore_read_enable;
  wire dp_sram_read_enable;
  wire [2:0] dp_sram_read_vector;
  wire pcore_read_wait;
  wire pcore_write_wait;
  wire [2:0] pcore_read_vector;
  wire [2:0] pcore_write_vector;
  wire pcore_write_stream;
  wire [1:0] pcore_write_stream_id;
  wire [1:0] pcore_read_data_flow;
  wire pcore_read_stream;
  wire [1:0] pcore_read_stream_id;
  wire [1:0] pcore_write_data_flow;
  wire [1:0] pcore_read_data_type;
  wire [1:0] pcore_read_data_model;
  wire [1:0] pcore_write_data_type;
  wire [1:0] pcore_write_data_model;
  wire [2:0] dp_pcore_read_vector;
  wire [2:0] dp_pcore_write_vector;
  wire dp_pcore_write_stream;
  wire [1:0] dp_pcore_write_stream_id;
  wire [2:0] ddr_read_vector;
  wire [2:0] ddr_write_vector;
  wire [1:0] dp_pcore_read_data_flow;
  wire dp_pcore_read_stream;
  wire [1:0] dp_pcore_write_data_flow;
  wire [1:0] dp_pcore_read_data_type;
  wire [1:0] dp_pcore_read_data_model;
  wire [1:0] dp_pcore_write_data_type;
  wire [1:0] dp_pcore_write_data_model;
  wire [1:0] pcore_read_scatter;
  wire [1:0] pcore_write_scatter;
  wire [1:0] pcore_read_scatter2;
  wire [1:0] pcore_write_scatter2;
  wire task_lockstep;
  wire [3:0] task_tid_mask;
  wire [27:0] task_iregister_auto;
  wire [1:0] task_data_model;
  wire [3:0] ddr_read_start;
  wire [3:0] ddr_read_end;
  wire ddr_tx_busy;
  wire n40_o;
  wire n41_o;
  wire [14:0] n43_o;
  wire n47_o;
  wire n48_o;
  wire n49_o;
  wire n50_o;
  wire n51_o;
  wire n52_o;
  wire n53_o;
  wire n54_o;
  wire n55_o;
  wire n56_o;
  wire n57_o;
  wire n58_o;
  wire n59_o;
  wire n60_o;
  wire n61_o;
  wire n62_o;
  wire [14:0] n63_o;
  wire n66_o;
  wire n67_o;
  wire n68_o;
  wire n70_o;
  wire n71_o;
  wire [1:0] n73_o;
  wire n74_o;
  wire n79_o;
  wire n81_o;
  wire n82_o;
  wire n83_o;
  wire [31:0] n86_o;
  wire n88_o;
  wire n89_o;
  wire n91_o;
  wire [23:0] n95_o;
  wire n98_o;
  wire n99_o;
  wire n101_o;
  wire [23:0] n105_o;
  wire n108_o;
  wire n109_o;
  wire n111_o;
  wire [23:0] n115_o;
  wire n117_o;
  wire n119_o;
  wire [23:0] n123_o;
  wire [47:0] n125_o;
  wire [47:0] n126_o;
  wire [47:0] n127_o;
  wire n130_o;
  wire n131_o;
  wire n132_o;
  wire [31:0] n135_o;
  wire n137_o;
  wire n138_o;
  wire n140_o;
  wire [23:0] n144_o;
  wire n147_o;
  wire n148_o;
  wire n150_o;
  wire [23:0] n154_o;
  wire n157_o;
  wire n158_o;
  wire n160_o;
  wire [23:0] n164_o;
  wire n166_o;
  wire n168_o;
  wire [23:0] n172_o;
  wire [47:0] n174_o;
  wire [47:0] n175_o;
  wire [47:0] n176_o;
  wire n179_o;
  wire n180_o;
  wire n182_o;
  wire [23:0] n184_o;
  wire n186_o;
  wire [23:0] n188_o;
  wire n190_o;
  wire [23:0] n192_o;
  wire [23:0] n194_o;
  wire [23:0] n195_o;
  wire [23:0] n196_o;
  wire [23:0] n197_o;
  wire axilite_i_n221;
  wire axilite_i_n222;
  wire axilite_i_n223;
  wire [31:0] axilite_i_n224;
  wire [1:0] axilite_i_n225;
  wire axilite_i_n226;
  wire axilite_i_n227;
  wire axilite_i_n228;
  wire [1:0] axilite_i_n229;
  wire [23:0] axilite_i_n230;
  wire [23:0] axilite_i_n231;
  wire axilite_i_n232;
  wire axilite_i_n233;
  wire [31:0] axilite_i_n234;
  wire axilite_i_axilite_arready_out;
  wire axilite_i_axilite_rvalid_out;
  wire axilite_i_axilite_rlast_out;
  wire [31:0] axilite_i_axilite_rdata_out;
  wire [1:0] axilite_i_axilite_rresp_out;
  wire axilite_i_axilite_awready_out;
  wire axilite_i_axilite_wready_out;
  wire axilite_i_axilite_bvalid_out;
  wire [1:0] axilite_i_axilite_bresp_out;
  wire [23:0] axilite_i_bus_waddr_out;
  wire [23:0] axilite_i_bus_raddr_out;
  wire axilite_i_bus_write_out;
  wire axilite_i_bus_read_out;
  wire [31:0] axilite_i_bus_writedata_out;
  wire sram_i_n263;
  wire sram_i_n264;
  wire [63:0] sram_i_n265;
  wire sram_i_dp_readdatavalid_out;
  wire sram_i_dp_readdatavalid_vm_out;
  wire [63:0] sram_i_dp_readdata_out;
  wire n272_o;
  wire n274_o;
  wire n275_o;
  wire n276_o;
  wire n278_o;
  wire n280_o;
  wire n281_o;
  wire n282_o;
  wire n286_o;
  wire n289_o;
  localparam n291_o = 1'b0;
  wire ddr_rx_i_n292;
  wire ddr_rx_i_n294;
  wire ddr_rx_i_n295;
  wire [63:0] ddr_rx_i_n296;
  wire ddr_rx_i_n297;
  wire [31:0] ddr_rx_i_n298;
  wire [2:0] ddr_rx_i_n299;
  wire ddr_rx_i_n300;
  wire ddr_rx_i_n301;
  wire [1:0] ddr_rx_i_n302;
  wire [3:0] ddr_rx_i_n303;
  wire ddr_rx_i_n304;
  wire ddr_rx_i_n305;
  wire [2:0] ddr_rx_i_n306;
  wire [3:0] ddr_rx_i_n307;
  wire [2:0] ddr_rx_i_n308;
  wire ddr_rx_i_read_data_ready_out;
  wire ddr_rx_i_read_fork_out;
  wire ddr_rx_i_read_data_valid_out;
  wire ddr_rx_i_read_data_valid_vm_out;
  wire [63:0] ddr_rx_i_read_data_out;
  wire ddr_rx_i_read_wait_request_out;
  wire [31:0] ddr_rx_i_ddr_araddr_out;
  wire [2:0] ddr_rx_i_ddr_arlen_out;
  wire ddr_rx_i_ddr_arvalid_out;
  wire ddr_rx_i_ddr_rready_out;
  wire [1:0] ddr_rx_i_ddr_arburst_out;
  wire [3:0] ddr_rx_i_ddr_arcache_out;
  wire ddr_rx_i_ddr_arid_out;
  wire ddr_rx_i_ddr_arlock_out;
  wire [2:0] ddr_rx_i_ddr_arprot_out;
  wire [3:0] ddr_rx_i_ddr_arqos_out;
  wire [2:0] ddr_rx_i_ddr_arsize_out;
  wire ddr_tx_i_n342;
  wire [31:0] ddr_tx_i_n343;
  wire [2:0] ddr_tx_i_n344;
  wire ddr_tx_i_n345;
  wire [31:0] ddr_tx_i_n346;
  wire ddr_tx_i_n347;
  wire [63:0] ddr_tx_i_n348;
  wire ddr_tx_i_n349;
  wire [7:0] ddr_tx_i_n350;
  wire [1:0] ddr_tx_i_n351;
  wire [3:0] ddr_tx_i_n352;
  wire ddr_tx_i_n353;
  wire ddr_tx_i_n354;
  wire [2:0] ddr_tx_i_n355;
  wire [3:0] ddr_tx_i_n356;
  wire [2:0] ddr_tx_i_n357;
  wire ddr_tx_i_n358;
  wire ddr_tx_i_n359;
  wire ddr_tx_i_write_wait_request_out;
  wire [31:0] ddr_tx_i_ddr_awaddr_out;
  wire [2:0] ddr_tx_i_ddr_awlen_out;
  wire ddr_tx_i_ddr_awvalid_out;
  wire [31:0] ddr_tx_i_ddr_waddr_out;
  wire ddr_tx_i_ddr_wvalid_out;
  wire [63:0] ddr_tx_i_ddr_wdata_out;
  wire ddr_tx_i_ddr_wlast_out;
  wire [7:0] ddr_tx_i_ddr_wbe_out;
  wire [1:0] ddr_tx_i_ddr_awburst_out;
  wire [3:0] ddr_tx_i_ddr_awcache_out;
  wire ddr_tx_i_ddr_awid_out;
  wire ddr_tx_i_ddr_awlock_out;
  wire [2:0] ddr_tx_i_ddr_awprot_out;
  wire [3:0] ddr_tx_i_ddr_awqos_out;
  wire [2:0] ddr_tx_i_ddr_awsize_out;
  wire ddr_tx_i_ddr_bready_out;
  wire ddr_tx_i_ddr_tx_busy_out;
  wire [11:0] n396_o;
  wire [11:0] n397_o;
  wire [31:0] dp_1_i_n398;
  wire dp_1_i_n399;
  wire dp_1_i_n400;
  wire dp_1_i_n401;
  wire [21:0] dp_1_i_n402;
  wire dp_1_i_n403;
  wire dp_1_i_n404;
  wire dp_1_i_n406;
  wire dp_1_i_n407;
  wire [1:0] dp_1_i_n408;
  wire dp_1_i_n409;
  wire [1:0] dp_1_i_n410;
  wire [2:0] dp_1_i_n411;
  wire [1:0] dp_1_i_n412;
  wire [1:0] dp_1_i_n415;
  wire [1:0] dp_1_i_n416;
  wire [21:0] dp_1_i_n417;
  wire dp_1_i_n418;
  wire dp_1_i_n419;
  wire dp_1_i_n420;
  wire [5:0] dp_1_i_n421;
  wire dp_1_i_n423;
  wire [1:0] dp_1_i_n424;
  wire [2:0] dp_1_i_n425;
  wire dp_1_i_n426;
  wire [1:0] dp_1_i_n427;
  wire [1:0] dp_1_i_n428;
  wire [63:0] dp_1_i_n429;
  wire [1:0] dp_1_i_n432;
  wire [1:0] dp_1_i_n433;
  wire [17:0] dp_1_i_n435;
  wire dp_1_i_n436;
  wire dp_1_i_n438;
  wire dp_1_i_n439;
  wire [2:0] dp_1_i_n440;
  wire [17:0] dp_1_i_n444;
  wire dp_1_i_n445;
  wire dp_1_i_n447;
  wire dp_1_i_n448;
  wire [2:0] dp_1_i_n449;
  wire [63:0] dp_1_i_n451;
  wire [31:0] dp_1_i_n455;
  wire dp_1_i_n457;
  wire dp_1_i_n458;
  wire [2:0] dp_1_i_n459;
  wire [3:0] dp_1_i_n461;
  wire [3:0] dp_1_i_n462;
  wire [4:0] dp_1_i_n463;
  wire [15:0] dp_1_i_n465;
  wire [31:0] dp_1_i_n466;
  wire dp_1_i_n468;
  wire [2:0] dp_1_i_n470;
  wire [3:0] dp_1_i_n472;
  wire [63:0] dp_1_i_n473;
  wire [4:0] dp_1_i_n474;
  wire [8:0] dp_1_i_n475;
  wire [4:0] dp_1_i_n476;
  wire [10:0] dp_1_i_n479;
  wire dp_1_i_n480;
  wire dp_1_i_n481;
  wire [4:0] dp_1_i_n482;
  wire dp_1_i_n483;
  wire [3:0] dp_1_i_n484;
  wire [27:0] dp_1_i_n485;
  wire [1:0] dp_1_i_n486;
  wire [1:0] dp_1_i_n487;
  wire [31:0] dp_1_i_bus_readdata_out;
  wire dp_1_i_bus_readdatavalid_out;
  wire dp_1_i_bus_writewait_out;
  wire dp_1_i_bus_readwait_out;
  wire [21:0] dp_1_i_readmaster1_addr_out;
  wire dp_1_i_readmaster1_fork_out;
  wire dp_1_i_readmaster1_addr_mode_out;
  wire dp_1_i_readmaster1_cs_out;
  wire dp_1_i_readmaster1_read_out;
  wire dp_1_i_readmaster1_read_vm_out;
  wire [1:0] dp_1_i_readmaster1_read_data_flow_out;
  wire dp_1_i_readmaster1_read_stream_out;
  wire [1:0] dp_1_i_readmaster1_read_stream_id_out;
  wire [2:0] dp_1_i_readmaster1_read_vector_out;
  wire [1:0] dp_1_i_readmaster1_read_scatter_out;
  wire [4:0] dp_1_i_readmaster1_burstlen_out;
  wire [1:0] dp_1_i_readmaster1_bus_id_out;
  wire [1:0] dp_1_i_readmaster1_data_type_out;
  wire [1:0] dp_1_i_readmaster1_data_model_out;
  wire [21:0] dp_1_i_writemaster1_addr_out;
  wire dp_1_i_writemaster1_fork_out;
  wire dp_1_i_writemaster1_addr_mode_out;
  wire dp_1_i_writemaster1_vm_out;
  wire [5:0] dp_1_i_writemaster1_mcast_out;
  wire dp_1_i_writemaster1_cs_out;
  wire dp_1_i_writemaster1_write_out;
  wire [1:0] dp_1_i_writemaster1_write_data_flow_out;
  wire [2:0] dp_1_i_writemaster1_write_vector_out;
  wire dp_1_i_writemaster1_write_stream_out;
  wire [1:0] dp_1_i_writemaster1_write_stream_id_out;
  wire [1:0] dp_1_i_writemaster1_write_scatter_out;
  wire [63:0] dp_1_i_writemaster1_writedata_out;
  wire [4:0] dp_1_i_writemaster1_burstlen_out;
  wire [1:0] dp_1_i_writemaster1_bus_id_out;
  wire [1:0] dp_1_i_writemaster1_data_type_out;
  wire [1:0] dp_1_i_writemaster1_data_model_out;
  wire dp_1_i_writemaster1_thread_out;
  wire [17:0] dp_1_i_readmaster2_addr_out;
  wire dp_1_i_readmaster2_fork_out;
  wire dp_1_i_readmaster2_cs_out;
  wire dp_1_i_readmaster2_read_out;
  wire dp_1_i_readmaster2_read_vm_out;
  wire [2:0] dp_1_i_readmaster2_read_vector_out;
  wire [1:0] dp_1_i_readmaster2_read_scatter_out;
  wire [4:0] dp_1_i_readmaster2_burstlen_out;
  wire [1:0] dp_1_i_readmaster2_bus_id_out;
  wire [17:0] dp_1_i_writemaster2_addr_out;
  wire dp_1_i_writemaster2_fork_out;
  wire dp_1_i_writemaster2_cs_out;
  wire dp_1_i_writemaster2_write_out;
  wire dp_1_i_writemaster2_vm_out;
  wire [2:0] dp_1_i_writemaster2_write_vector_out;
  wire [1:0] dp_1_i_writemaster2_write_scatter_out;
  wire [63:0] dp_1_i_writemaster2_writedata_out;
  wire [4:0] dp_1_i_writemaster2_burstlen_out;
  wire [1:0] dp_1_i_writemaster2_bus_id_out;
  wire dp_1_i_writemaster2_thread_out;
  wire [31:0] dp_1_i_readmaster3_addr_out;
  wire dp_1_i_readmaster3_cs_out;
  wire dp_1_i_readmaster3_read_out;
  wire dp_1_i_readmaster3_read_vm_out;
  wire [2:0] dp_1_i_readmaster3_read_vector_out;
  wire [1:0] dp_1_i_readmaster3_read_scatter_out;
  wire [3:0] dp_1_i_readmaster3_read_start_out;
  wire [3:0] dp_1_i_readmaster3_read_end_out;
  wire [4:0] dp_1_i_readmaster3_burstlen_out;
  wire [1:0] dp_1_i_readmaster3_bus_id_out;
  wire [15:0] dp_1_i_readmaster3_filler_data_out;
  wire [31:0] dp_1_i_writemaster3_addr_out;
  wire dp_1_i_writemaster3_cs_out;
  wire dp_1_i_writemaster3_write_out;
  wire dp_1_i_writemaster3_vm_out;
  wire [2:0] dp_1_i_writemaster3_write_vector_out;
  wire [1:0] dp_1_i_writemaster3_write_scatter_out;
  wire [3:0] dp_1_i_writemaster3_write_end_out;
  wire [63:0] dp_1_i_writemaster3_writedata_out;
  wire [4:0] dp_1_i_writemaster3_burstlen_out;
  wire [8:0] dp_1_i_writemaster3_burstlen2_out;
  wire [4:0] dp_1_i_writemaster3_burstlen3_out;
  wire [1:0] dp_1_i_writemaster3_bus_id_out;
  wire dp_1_i_writemaster3_thread_out;
  wire [15:0] dp_1_i_writemaster3_filler_data_out;
  wire [10:0] dp_1_i_task_start_addr_out;
  wire dp_1_i_task_out;
  wire dp_1_i_task_vm_out;
  wire [4:0] dp_1_i_task_pcore_out;
  wire dp_1_i_task_lockstep_out;
  wire [3:0] dp_1_i_task_tid_mask_out;
  wire [27:0] dp_1_i_task_iregister_auto_out;
  wire [1:0] dp_1_i_task_data_model_out;
  wire [1:0] dp_1_i_task_busy_out;
  wire dp_1_i_indication_avail_out;
  wire core_i_n646;
  wire core_i_n647;
  wire core_i_n648;
  wire core_i_n649;
  wire [63:0] core_i_n650;
  wire core_i_n651;
  wire [1:0] core_i_n652;
  wire core_i_n653;
  wire core_i_dp_write_wait_out;
  wire core_i_dp_read_wait_out;
  wire core_i_dp_readdatavalid_out;
  wire core_i_dp_read_gen_valid_out;
  wire [63:0] core_i_dp_readdata_out;
  wire core_i_dp_readdata_vm_out;
  wire [1:0] core_i_busy_out;
  wire core_i_ready_out;
  wire [71:0] n670_o;
  wire [47:0] n671_o;
  reg [47:0] n672_q;
  wire [47:0] n673_o;
  reg [47:0] n674_q;
  wire [23:0] n675_o;
  reg [23:0] n676_q;
  wire [23:0] n678_o;
  wire [23:0] n679_o;
  wire [23:0] n680_o;
  wire n681_o;
  wire n682_o;
  wire [23:0] n683_o;
  wire [23:0] n684_o;
  wire [23:0] n685_o;
  wire [23:0] n686_o;
  wire [47:0] n687_o;
  wire [23:0] n688_o;
  wire [23:0] n689_o;
  wire [23:0] n690_o;
  wire n691_o;
  wire n692_o;
  wire [23:0] n693_o;
  wire [23:0] n694_o;
  wire [23:0] n695_o;
  wire [23:0] n696_o;
  wire [47:0] n697_o;
  wire [23:0] n698_o;
  wire [23:0] n699_o;
  wire [23:0] n700_o;
  wire n701_o;
  wire n702_o;
  wire [23:0] n703_o;
  wire [23:0] n704_o;
  wire [23:0] n705_o;
  wire [23:0] n706_o;
  wire [47:0] n707_o;
  wire [23:0] n708_o;
  wire [23:0] n709_o;
  wire [23:0] n710_o;
  wire n711_o;
  wire n712_o;
  wire [23:0] n713_o;
  wire [23:0] n714_o;
  wire [23:0] n715_o;
  wire [23:0] n716_o;
  wire [47:0] n717_o;
  wire [23:0] n718_o;
  wire [23:0] n719_o;
  wire [23:0] n720_o;
  wire n721_o;
  wire n722_o;
  wire [23:0] n723_o;
  wire [23:0] n724_o;
  wire [23:0] n725_o;
  wire [23:0] n726_o;
  wire [47:0] n727_o;
  wire [23:0] n728_o;
  wire [23:0] n729_o;
  wire [23:0] n730_o;
  wire n731_o;
  wire n732_o;
  wire [23:0] n733_o;
  wire [23:0] n734_o;
  wire [23:0] n735_o;
  wire [23:0] n736_o;
  wire [47:0] n737_o;
  wire [23:0] n738_o;
  wire [23:0] n739_o;
  wire [23:0] n740_o;
  wire n741_o;
  wire n742_o;
  wire [23:0] n743_o;
  wire [23:0] n744_o;
  wire [23:0] n745_o;
  wire [23:0] n746_o;
  wire [47:0] n747_o;
  wire [23:0] n748_o;
  wire [23:0] n749_o;
  wire [23:0] n750_o;
  wire n751_o;
  wire n752_o;
  wire [23:0] n753_o;
  wire [23:0] n754_o;
  wire [23:0] n755_o;
  wire [23:0] n756_o;
  wire [47:0] n757_o;
  assign axi_araddr_out = ddr_rx_i_n298;
  assign axi_arlen_out = ddr_rx_i_n299;
  assign axi_arvalid_out = ddr_rx_i_n300;
  assign axi_rready_out = ddr_rx_i_n301;
  assign axi_arburst_out = ddr_rx_i_n302;
  assign axi_arcache_out = ddr_rx_i_n303;
  assign axi_arid_out = ddr_rx_i_n304;
  assign axi_arlock_out = ddr_rx_i_n305;
  assign axi_arprot_out = ddr_rx_i_n306;
  assign axi_arqos_out = ddr_rx_i_n307;
  assign axi_arsize_out = ddr_rx_i_n308;
  assign axi_awaddr_out = ddr_tx_i_n343;
  assign axi_awlen_out = ddr_tx_i_n344;
  assign axi_awvalid_out = ddr_tx_i_n345;
  assign axi_waddr_out = ddr_tx_i_n346;
  assign axi_wvalid_out = ddr_tx_i_n347;
  assign axi_wdata_out = ddr_tx_i_n348;
  assign axi_wlast_out = ddr_tx_i_n349;
  assign axi_wbe_out = ddr_tx_i_n350;
  assign axi_awburst_out = ddr_tx_i_n351;
  assign axi_awcache_out = ddr_tx_i_n352;
  assign axi_awid_out = ddr_tx_i_n353;
  assign axi_awlock_out = ddr_tx_i_n354;
  assign axi_awprot_out = ddr_tx_i_n355;
  assign axi_awqos_out = ddr_tx_i_n356;
  assign axi_awsize_out = ddr_tx_i_n357;
  assign axi_bready_out = ddr_tx_i_n358;
  assign axilite_arready_out = axilite_i_n221;
  assign axilite_rvalid_out = axilite_i_n222;
  assign axilite_rlast_out = axilite_i_n223;
  assign axilite_rdata_out = axilite_i_n224;
  assign axilite_rresp_out = axilite_i_n225;
  assign axilite_awready_out = axilite_i_n226;
  assign axilite_wready_out = axilite_i_n227;
  assign axilite_bvalid_out = axilite_i_n228;
  assign axilite_bresp_out = axilite_i_n229;
  /* ../../HW/src/top/ztachip.vhd:100:8  */
  assign host_waddr = axilite_i_n230; // (signal)
  /* ../../HW/src/top/ztachip.vhd:101:8  */
  assign host_raddr = axilite_i_n231; // (signal)
  /* ../../HW/src/top/ztachip.vhd:102:8  */
  assign host_wren = axilite_i_n232; // (signal)
  /* ../../HW/src/top/ztachip.vhd:103:8  */
  assign host_rden = axilite_i_n233; // (signal)
  /* ../../HW/src/top/ztachip.vhd:104:8  */
  assign host_writedata = axilite_i_n234; // (signal)
  /* ../../HW/src/top/ztachip.vhd:105:8  */
  assign host_readdata = dp_1_i_n398; // (signal)
  /* ../../HW/src/top/ztachip.vhd:106:8  */
  assign host_readdatavalid = dp_1_i_n399; // (signal)
  /* ../../HW/src/top/ztachip.vhd:107:8  */
  assign host_writewait = dp_1_i_n400; // (signal)
  /* ../../HW/src/top/ztachip.vhd:108:8  */
  assign host_readwait = dp_1_i_n401; // (signal)
  /* ../../HW/src/top/ztachip.vhd:112:8  */
  assign pcore_busy = dp_1_i_n487; // (signal)
  /* ../../HW/src/top/ztachip.vhd:113:8  */
  assign busy = core_i_n652; // (signal)
  /* ../../HW/src/top/ztachip.vhd:114:8  */
  assign pcore_read_busy = n53_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:115:8  */
  assign pcore_write_busy = n60_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:116:8  */
  assign ready = core_i_n653; // (signal)
  /* ../../HW/src/top/ztachip.vhd:120:8  */
  assign pcore_read_addr = dp_pcore_read_addr; // (signal)
  /* ../../HW/src/top/ztachip.vhd:121:8  */
  assign pcore_read_fork = dp_pcore_read_fork; // (signal)
  /* ../../HW/src/top/ztachip.vhd:122:8  */
  assign pcore_read_addr_mode = dp_pcore_read_addr_mode; // (signal)
  /* ../../HW/src/top/ztachip.vhd:123:8  */
  assign pcore_read_enable = n41_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:124:8  */
  assign pcore_read_gen_valid = 1'b1; // (signal)
  /* ../../HW/src/top/ztachip.vhd:125:8  */
  assign pcore_read_data = core_i_n650; // (signal)
  /* ../../HW/src/top/ztachip.vhd:126:8  */
  assign pcore_readdata_vm = core_i_n651; // (signal)
  /* ../../HW/src/top/ztachip.vhd:127:8  */
  assign pcore_read_data_valid = core_i_n648; // (signal)
  /* ../../HW/src/top/ztachip.vhd:128:8  */
  assign pcore_read_data_valid2 = n74_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:129:8  */
  assign pcore_read_gen_valid2 = core_i_n649; // (signal)
  /* ../../HW/src/top/ztachip.vhd:133:8  */
  assign pcore_write_addr = dp_pcore_write_addr; // (signal)
  /* ../../HW/src/top/ztachip.vhd:134:8  */
  assign pcore_write_fork = dp_pcore_write_fork; // (signal)
  /* ../../HW/src/top/ztachip.vhd:135:8  */
  assign pcore_write_addr_mode = dp_1_i_n419; // (signal)
  /* ../../HW/src/top/ztachip.vhd:136:8  */
  assign pcore_mcast = dp_1_i_n421; // (signal)
  /* ../../HW/src/top/ztachip.vhd:137:8  */
  assign pcore_write_enable = n71_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:138:8  */
  assign pcore_write_gen_valid = 1'b1; // (signal)
  /* ../../HW/src/top/ztachip.vhd:139:8  */
  assign pcore_write_data = dp_pcore_write_data; // (signal)
  /* ../../HW/src/top/ztachip.vhd:143:8  */
  assign sram_read_addr = n43_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:144:8  */
  assign sram_read_fork = dp_sram_read_fork; // (signal)
  /* ../../HW/src/top/ztachip.vhd:145:8  */
  assign sram_read_enable = dp_sram_read_enable; // (signal)
  /* ../../HW/src/top/ztachip.vhd:146:8  */
  assign sram_read_vector = dp_sram_read_vector; // (signal)
  /* ../../HW/src/top/ztachip.vhd:147:8  */
  assign sram_read_gen_valid = 1'b1; // (signal)
  /* ../../HW/src/top/ztachip.vhd:148:8  */
  assign sram_read_data = sram_i_n265; // (signal)
  /* ../../HW/src/top/ztachip.vhd:149:8  */
  assign sram_read_data_valid = sram_i_n263; // (signal)
  /* ../../HW/src/top/ztachip.vhd:150:8  */
  assign sram_readdata_vm = sram_i_n264; // (signal)
  /* ../../HW/src/top/ztachip.vhd:151:8  */
  assign sram_read_vm = dp_1_i_n439; // (signal)
  /* ../../HW/src/top/ztachip.vhd:155:8  */
  assign sram_write_addr = n63_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:156:8  */
  assign sram_write_fork = dp_sram_write_fork; // (signal)
  /* ../../HW/src/top/ztachip.vhd:157:8  */
  assign sram_write_enable = n68_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:158:8  */
  assign sram_write_vector = dp_sram_write_vector; // (signal)
  /* ../../HW/src/top/ztachip.vhd:159:8  */
  assign sram_write_data = dp_sram_write_data; // (signal)
  /* ../../HW/src/top/ztachip.vhd:163:8  */
  assign ddr_read_addr = dp_1_i_n455; // (signal)
  /* ../../HW/src/top/ztachip.vhd:164:8  */
  assign ddr_read_enable = dp_1_i_n457; // (signal)
  /* ../../HW/src/top/ztachip.vhd:165:8  */
  assign ddr_read_enable_2 = n276_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:166:8  */
  assign ddr_read_wait = ddr_rx_i_n297; // (signal)
  /* ../../HW/src/top/ztachip.vhd:167:8  */
  assign ddr_read_wait_2 = n272_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:168:8  */
  assign ddr_read_data = ddr_rx_i_n296; // (signal)
  /* ../../HW/src/top/ztachip.vhd:169:8  */
  assign ddr_read_data_valid = ddr_rx_i_n294; // (signal)
  /* ../../HW/src/top/ztachip.vhd:170:8  */
  assign ddr_read_burstlen = dp_1_i_n463; // (signal)
  /* ../../HW/src/top/ztachip.vhd:171:8  */
  assign ddr_read_filler_data = dp_1_i_n465; // (signal)
  /* ../../HW/src/top/ztachip.vhd:175:8  */
  assign ddr_write_addr = dp_1_i_n466; // (signal)
  /* ../../HW/src/top/ztachip.vhd:176:8  */
  assign ddr_write_enable = dp_1_i_n468; // (signal)
  /* ../../HW/src/top/ztachip.vhd:177:8  */
  assign ddr_write_enable_2 = n282_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:178:8  */
  assign ddr_write_wait = ddr_tx_i_n342; // (signal)
  /* ../../HW/src/top/ztachip.vhd:179:8  */
  assign ddr_write_wait_2 = n278_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:180:8  */
  assign ddr_write_data = dp_1_i_n473; // (signal)
  /* ../../HW/src/top/ztachip.vhd:181:8  */
  assign ddr_write_burstlen = dp_1_i_n474; // (signal)
  /* ../../HW/src/top/ztachip.vhd:182:8  */
  assign ddr_write_burstlen2 = dp_1_i_n475; // (signal)
  /* ../../HW/src/top/ztachip.vhd:183:8  */
  assign ddr_write_burstlen3 = dp_1_i_n476; // (signal)
  /* ../../HW/src/top/ztachip.vhd:185:8  */
  assign ddr_data_ready = ddr_rx_i_n292; // (signal)
  /* ../../HW/src/top/ztachip.vhd:186:8  */
  assign ddr_data_wait = n289_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:187:8  */
  assign ddr_write_end = dp_1_i_n472; // (signal)
  /* ../../HW/src/top/ztachip.vhd:188:8  */
  assign ddr_read_vm = dp_1_i_n458; // (signal)
  /* ../../HW/src/top/ztachip.vhd:189:8  */
  assign ddr_readdata_vm = ddr_rx_i_n295; // (signal)
  /* ../../HW/src/top/ztachip.vhd:193:8  */
  assign task_start_addr = dp_1_i_n479; // (signal)
  /* ../../HW/src/top/ztachip.vhd:194:8  */
  assign \task  = dp_1_i_n480; // (signal)
  /* ../../HW/src/top/ztachip.vhd:195:8  */
  assign task_vm = dp_1_i_n481; // (signal)
  /* ../../HW/src/top/ztachip.vhd:196:8  */
  assign task_pcore = dp_1_i_n482; // (signal)
  /* ../../HW/src/top/ztachip.vhd:198:8  */
  assign bar = n670_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:202:8  */
  assign pcore_write_counter_r = n672_q; // (signal)
  /* ../../HW/src/top/ztachip.vhd:203:8  */
  assign sram_write_counter_r = n674_q; // (signal)
  /* ../../HW/src/top/ztachip.vhd:204:8  */
  assign ddr_write_counter_r = n676_q; // (signal)
  /* ../../HW/src/top/ztachip.vhd:206:8  */
  assign dp_sram_read_fork = dp_1_i_n436; // (signal)
  /* ../../HW/src/top/ztachip.vhd:207:8  */
  assign dp_sram_read_wait = 1'b0; // (signal)
  /* ../../HW/src/top/ztachip.vhd:208:8  */
  assign dp_sram_write_fork = dp_1_i_n445; // (signal)
  /* ../../HW/src/top/ztachip.vhd:209:8  */
  assign dp_sram_write_wait = 1'b0; // (signal)
  /* ../../HW/src/top/ztachip.vhd:210:8  */
  assign dp_sram_write_enable = dp_1_i_n447; // (signal)
  /* ../../HW/src/top/ztachip.vhd:211:8  */
  assign dp_sram_write_vector = dp_1_i_n449; // (signal)
  /* ../../HW/src/top/ztachip.vhd:212:8  */
  assign dp_sram_write_addr = dp_1_i_n444; // (signal)
  /* ../../HW/src/top/ztachip.vhd:213:8  */
  assign dp_sram_write_data = dp_1_i_n451; // (signal)
  /* ../../HW/src/top/ztachip.vhd:214:8  */
  assign dp_sram_write_page = n73_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:215:8  */
  assign dp_sram_write_vm = dp_1_i_n448; // (signal)
  /* ../../HW/src/top/ztachip.vhd:217:8  */
  assign dp_pcore_read_wait = n61_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:218:8  */
  assign dp_pcore_write_wait = n62_o; // (signal)
  /* ../../HW/src/top/ztachip.vhd:219:8  */
  assign dp_pcore_write_addr = dp_1_i_n417; // (signal)
  /* ../../HW/src/top/ztachip.vhd:220:8  */
  assign dp_pcore_write_fork = dp_1_i_n418; // (signal)
  /* ../../HW/src/top/ztachip.vhd:221:8  */
  assign dp_pcore_write_data = dp_1_i_n429; // (signal)
  /* ../../HW/src/top/ztachip.vhd:222:8  */
  assign dp_pcore_write_enable = dp_1_i_n423; // (signal)
  /* ../../HW/src/top/ztachip.vhd:223:8  */
  assign dp_pcore_write_vm = dp_1_i_n420; // (signal)
  /* ../../HW/src/top/ztachip.vhd:224:8  */
  assign dp_pcore_read_vm = dp_1_i_n407; // (signal)
  /* ../../HW/src/top/ztachip.vhd:226:8  */
  assign dp_pcore_read_addr = dp_1_i_n402; // (signal)
  /* ../../HW/src/top/ztachip.vhd:227:8  */
  assign dp_pcore_read_fork = dp_1_i_n403; // (signal)
  /* ../../HW/src/top/ztachip.vhd:228:8  */
  assign dp_pcore_read_addr_mode = dp_1_i_n404; // (signal)
  /* ../../HW/src/top/ztachip.vhd:229:8  */
  assign dp_sram_read_addr = dp_1_i_n435; // (signal)
  /* ../../HW/src/top/ztachip.vhd:230:8  */
  assign dp_pcore_read_enable = dp_1_i_n406; // (signal)
  /* ../../HW/src/top/ztachip.vhd:231:8  */
  assign dp_sram_read_enable = dp_1_i_n438; // (signal)
  /* ../../HW/src/top/ztachip.vhd:232:8  */
  assign dp_sram_read_vector = dp_1_i_n440; // (signal)
  /* ../../HW/src/top/ztachip.vhd:234:8  */
  assign pcore_read_wait = core_i_n647; // (signal)
  /* ../../HW/src/top/ztachip.vhd:235:8  */
  assign pcore_write_wait = core_i_n646; // (signal)
  /* ../../HW/src/top/ztachip.vhd:237:8  */
  assign pcore_read_vector = dp_pcore_read_vector; // (signal)
  /* ../../HW/src/top/ztachip.vhd:238:8  */
  assign pcore_write_vector = dp_pcore_write_vector; // (signal)
  /* ../../HW/src/top/ztachip.vhd:239:8  */
  assign pcore_write_stream = dp_pcore_write_stream; // (signal)
  /* ../../HW/src/top/ztachip.vhd:240:8  */
  assign pcore_write_stream_id = dp_pcore_write_stream_id; // (signal)
  /* ../../HW/src/top/ztachip.vhd:241:8  */
  assign pcore_read_data_flow = dp_pcore_read_data_flow; // (signal)
  /* ../../HW/src/top/ztachip.vhd:242:8  */
  assign pcore_read_stream = dp_pcore_read_stream; // (signal)
  /* ../../HW/src/top/ztachip.vhd:243:8  */
  assign pcore_read_stream_id = dp_1_i_n410; // (signal)
  /* ../../HW/src/top/ztachip.vhd:244:8  */
  assign pcore_write_data_flow = dp_pcore_write_data_flow; // (signal)
  /* ../../HW/src/top/ztachip.vhd:245:8  */
  assign pcore_read_data_type = dp_pcore_read_data_type; // (signal)
  /* ../../HW/src/top/ztachip.vhd:246:8  */
  assign pcore_read_data_model = dp_pcore_read_data_model; // (signal)
  /* ../../HW/src/top/ztachip.vhd:247:8  */
  assign pcore_write_data_type = dp_pcore_write_data_type; // (signal)
  /* ../../HW/src/top/ztachip.vhd:248:8  */
  assign pcore_write_data_model = dp_pcore_write_data_model; // (signal)
  /* ../../HW/src/top/ztachip.vhd:249:8  */
  assign dp_pcore_read_vector = dp_1_i_n411; // (signal)
  /* ../../HW/src/top/ztachip.vhd:250:8  */
  assign dp_pcore_write_vector = dp_1_i_n425; // (signal)
  /* ../../HW/src/top/ztachip.vhd:251:8  */
  assign dp_pcore_write_stream = dp_1_i_n426; // (signal)
  /* ../../HW/src/top/ztachip.vhd:252:8  */
  assign dp_pcore_write_stream_id = dp_1_i_n427; // (signal)
  /* ../../HW/src/top/ztachip.vhd:253:8  */
  assign ddr_read_vector = dp_1_i_n459; // (signal)
  /* ../../HW/src/top/ztachip.vhd:254:8  */
  assign ddr_write_vector = dp_1_i_n470; // (signal)
  /* ../../HW/src/top/ztachip.vhd:255:8  */
  assign dp_pcore_read_data_flow = dp_1_i_n408; // (signal)
  /* ../../HW/src/top/ztachip.vhd:256:8  */
  assign dp_pcore_read_stream = dp_1_i_n409; // (signal)
  /* ../../HW/src/top/ztachip.vhd:257:8  */
  assign dp_pcore_write_data_flow = dp_1_i_n424; // (signal)
  /* ../../HW/src/top/ztachip.vhd:258:8  */
  assign dp_pcore_read_data_type = dp_1_i_n415; // (signal)
  /* ../../HW/src/top/ztachip.vhd:259:8  */
  assign dp_pcore_read_data_model = dp_1_i_n416; // (signal)
  /* ../../HW/src/top/ztachip.vhd:260:8  */
  assign dp_pcore_write_data_type = dp_1_i_n432; // (signal)
  /* ../../HW/src/top/ztachip.vhd:261:8  */
  assign dp_pcore_write_data_model = dp_1_i_n433; // (signal)
  /* ../../HW/src/top/ztachip.vhd:263:8  */
  assign pcore_read_scatter = dp_1_i_n412; // (signal)
  /* ../../HW/src/top/ztachip.vhd:264:8  */
  assign pcore_write_scatter = dp_1_i_n428; // (signal)
  /* ../../HW/src/top/ztachip.vhd:266:8  */
  assign pcore_read_scatter2 = pcore_read_scatter; // (signal)
  /* ../../HW/src/top/ztachip.vhd:267:8  */
  assign pcore_write_scatter2 = pcore_write_scatter; // (signal)
  /* ../../HW/src/top/ztachip.vhd:269:8  */
  assign task_lockstep = dp_1_i_n483; // (signal)
  /* ../../HW/src/top/ztachip.vhd:270:8  */
  assign task_tid_mask = dp_1_i_n484; // (signal)
  /* ../../HW/src/top/ztachip.vhd:271:8  */
  assign task_iregister_auto = dp_1_i_n485; // (signal)
  /* ../../HW/src/top/ztachip.vhd:272:8  */
  assign task_data_model = dp_1_i_n486; // (signal)
  /* ../../HW/src/top/ztachip.vhd:274:8  */
  assign ddr_read_start = dp_1_i_n461; // (signal)
  /* ../../HW/src/top/ztachip.vhd:275:8  */
  assign ddr_read_end = dp_1_i_n462; // (signal)
  /* ../../HW/src/top/ztachip.vhd:278:8  */
  assign ddr_tx_busy = ddr_tx_i_n359; // (signal)
  /* ../../HW/src/top/ztachip.vhd:291:48  */
  assign n40_o = ~pcore_read_busy;
  /* ../../HW/src/top/ztachip.vhd:291:43  */
  assign n41_o = dp_pcore_read_enable & n40_o;
  /* ../../HW/src/top/ztachip.vhd:303:36  */
  assign n43_o = dp_sram_read_addr[14:0];
  /* ../../HW/src/top/ztachip.vhd:316:48  */
  assign n47_o = ~dp_pcore_read_vm;
  /* ../../HW/src/top/ztachip.vhd:316:84  */
  assign n48_o = pcore_busy[0];
  /* ../../HW/src/top/ztachip.vhd:316:70  */
  assign n49_o = n47_o & n48_o;
  /* ../../HW/src/top/ztachip.vhd:316:124  */
  assign n50_o = pcore_busy[1];
  /* ../../HW/src/top/ztachip.vhd:316:110  */
  assign n51_o = dp_pcore_read_vm & n50_o;
  /* ../../HW/src/top/ztachip.vhd:316:89  */
  assign n52_o = n49_o | n51_o;
  /* ../../HW/src/top/ztachip.vhd:316:41  */
  assign n53_o = dp_pcore_read_enable & n52_o;
  /* ../../HW/src/top/ztachip.vhd:317:50  */
  assign n54_o = ~dp_pcore_write_vm;
  /* ../../HW/src/top/ztachip.vhd:317:87  */
  assign n55_o = pcore_busy[0];
  /* ../../HW/src/top/ztachip.vhd:317:73  */
  assign n56_o = n54_o & n55_o;
  /* ../../HW/src/top/ztachip.vhd:317:128  */
  assign n57_o = pcore_busy[1];
  /* ../../HW/src/top/ztachip.vhd:317:114  */
  assign n58_o = dp_pcore_write_vm & n57_o;
  /* ../../HW/src/top/ztachip.vhd:317:92  */
  assign n59_o = n56_o | n58_o;
  /* ../../HW/src/top/ztachip.vhd:317:43  */
  assign n60_o = dp_pcore_write_enable & n59_o;
  /* ../../HW/src/top/ztachip.vhd:319:39  */
  assign n61_o = pcore_read_busy | pcore_read_wait;
  /* ../../HW/src/top/ztachip.vhd:320:41  */
  assign n62_o = pcore_write_busy | pcore_write_wait;
  /* ../../HW/src/top/ztachip.vhd:325:38  */
  assign n63_o = dp_sram_write_addr[14:0];
  /* ../../HW/src/top/ztachip.vhd:326:79  */
  assign n66_o = dp_sram_write_page == 2'b00;
  /* ../../HW/src/top/ztachip.vhd:326:57  */
  assign n67_o = n66_o & dp_sram_write_enable;
  /* ../../HW/src/top/ztachip.vhd:326:26  */
  assign n68_o = n67_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ztachip.vhd:336:50  */
  assign n70_o = ~pcore_write_busy;
  /* ../../HW/src/top/ztachip.vhd:336:45  */
  assign n71_o = dp_pcore_write_enable & n70_o;
  /* ../../HW/src/top/ztachip.vhd:348:41  */
  assign n73_o = dp_sram_write_addr[17:16];
  /* ../../HW/src/top/ztachip.vhd:352:49  */
  assign n74_o = pcore_read_data_valid & pcore_read_gen_valid2;
  /* ../../HW/src/top/ztachip.vhd:362:17  */
  assign n79_o = ~reset_in;
  /* ../../HW/src/top/ztachip.vhd:368:65  */
  assign n81_o = ~dp_pcore_write_wait;
  /* ../../HW/src/top/ztachip.vhd:368:42  */
  assign n82_o = n81_o & dp_pcore_write_enable;
  /* ../../HW/src/top/ztachip.vhd:369:37  */
  assign n83_o = ~dp_pcore_write_vm;
  /* ../../HW/src/top/ztachip.vhd:369:17  */
  assign n86_o = n83_o ? 32'b00000000000000000000000000000000 : 32'b00000000000000000000000000000001;
  /* ../../HW/src/top/ztachip.vhd:374:41  */
  assign n88_o = dp_pcore_write_vector == 3'b001;
  /* ../../HW/src/top/ztachip.vhd:375:42  */
  assign n89_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:375:73  */
  assign n91_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:375:78  */
  assign n95_o = n680_o + 24'b000000000000000000000010;
  /* ../../HW/src/top/ztachip.vhd:376:44  */
  assign n98_o = dp_pcore_write_vector == 3'b011;
  /* ../../HW/src/top/ztachip.vhd:377:42  */
  assign n99_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:377:73  */
  assign n101_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:377:78  */
  assign n105_o = n690_o + 24'b000000000000000000000100;
  /* ../../HW/src/top/ztachip.vhd:378:44  */
  assign n108_o = dp_pcore_write_vector == 3'b111;
  /* ../../HW/src/top/ztachip.vhd:379:42  */
  assign n109_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:379:73  */
  assign n111_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:379:78  */
  assign n115_o = n700_o + 24'b000000000000000000001000;
  /* ../../HW/src/top/ztachip.vhd:381:42  */
  assign n117_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:381:73  */
  assign n119_o = n86_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:381:78  */
  assign n123_o = n710_o + 24'b000000000000000000000001;
  /* ../../HW/src/top/ztachip.vhd:378:17  */
  assign n125_o = n108_o ? n707_o : n717_o;
  /* ../../HW/src/top/ztachip.vhd:376:17  */
  assign n126_o = n98_o ? n697_o : n125_o;
  /* ../../HW/src/top/ztachip.vhd:374:17  */
  assign n127_o = n88_o ? n687_o : n126_o;
  /* ../../HW/src/top/ztachip.vhd:384:63  */
  assign n130_o = ~dp_sram_write_wait;
  /* ../../HW/src/top/ztachip.vhd:384:41  */
  assign n131_o = n130_o & dp_sram_write_enable;
  /* ../../HW/src/top/ztachip.vhd:385:36  */
  assign n132_o = ~dp_sram_write_vm;
  /* ../../HW/src/top/ztachip.vhd:385:17  */
  assign n135_o = n132_o ? 32'b00000000000000000000000000000000 : 32'b00000000000000000000000000000001;
  /* ../../HW/src/top/ztachip.vhd:390:40  */
  assign n137_o = dp_sram_write_vector == 3'b001;
  /* ../../HW/src/top/ztachip.vhd:391:41  */
  assign n138_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:391:76  */
  assign n140_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:391:86  */
  assign n144_o = n720_o + 24'b000000000000000000000010;
  /* ../../HW/src/top/ztachip.vhd:392:43  */
  assign n147_o = dp_sram_write_vector == 3'b011;
  /* ../../HW/src/top/ztachip.vhd:393:41  */
  assign n148_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:393:76  */
  assign n150_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:393:86  */
  assign n154_o = n730_o + 24'b000000000000000000000100;
  /* ../../HW/src/top/ztachip.vhd:394:43  */
  assign n157_o = dp_sram_write_vector == 3'b111;
  /* ../../HW/src/top/ztachip.vhd:395:41  */
  assign n158_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:395:76  */
  assign n160_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:395:86  */
  assign n164_o = n740_o + 24'b000000000000000000001000;
  /* ../../HW/src/top/ztachip.vhd:397:41  */
  assign n166_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:397:76  */
  assign n168_o = n135_o[0];  // trunc
  /* ../../HW/src/top/ztachip.vhd:397:86  */
  assign n172_o = n750_o + 24'b000000000000000000000001;
  /* ../../HW/src/top/ztachip.vhd:394:17  */
  assign n174_o = n157_o ? n747_o : n757_o;
  /* ../../HW/src/top/ztachip.vhd:392:17  */
  assign n175_o = n147_o ? n737_o : n174_o;
  /* ../../HW/src/top/ztachip.vhd:390:17  */
  assign n176_o = n137_o ? n727_o : n175_o;
  /* ../../HW/src/top/ztachip.vhd:400:57  */
  assign n179_o = ~ddr_write_wait_2;
  /* ../../HW/src/top/ztachip.vhd:400:37  */
  assign n180_o = n179_o & ddr_write_enable;
  /* ../../HW/src/top/ztachip.vhd:401:36  */
  assign n182_o = ddr_write_vector == 3'b001;
  /* ../../HW/src/top/ztachip.vhd:402:62  */
  assign n184_o = ddr_write_counter_r + 24'b000000000000000000000010;
  /* ../../HW/src/top/ztachip.vhd:403:39  */
  assign n186_o = ddr_write_vector == 3'b011;
  /* ../../HW/src/top/ztachip.vhd:404:62  */
  assign n188_o = ddr_write_counter_r + 24'b000000000000000000000100;
  /* ../../HW/src/top/ztachip.vhd:405:39  */
  assign n190_o = ddr_write_vector == 3'b111;
  /* ../../HW/src/top/ztachip.vhd:406:62  */
  assign n192_o = ddr_write_counter_r + 24'b000000000000000000001000;
  /* ../../HW/src/top/ztachip.vhd:408:62  */
  assign n194_o = ddr_write_counter_r + 24'b000000000000000000000001;
  /* ../../HW/src/top/ztachip.vhd:405:17  */
  assign n195_o = n190_o ? n192_o : n194_o;
  /* ../../HW/src/top/ztachip.vhd:403:17  */
  assign n196_o = n186_o ? n188_o : n195_o;
  /* ../../HW/src/top/ztachip.vhd:401:17  */
  assign n197_o = n182_o ? n184_o : n196_o;
  /* ../../HW/src/top/ztachip.vhd:426:30  */
  assign axilite_i_n221 = axilite_i_axilite_arready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:427:29  */
  assign axilite_i_n222 = axilite_i_axilite_rvalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:428:28  */
  assign axilite_i_n223 = axilite_i_axilite_rlast_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:429:28  */
  assign axilite_i_n224 = axilite_i_axilite_rdata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:431:28  */
  assign axilite_i_n225 = axilite_i_axilite_rresp_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:437:30  */
  assign axilite_i_n226 = axilite_i_axilite_awready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:438:29  */
  assign axilite_i_n227 = axilite_i_axilite_wready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:439:29  */
  assign axilite_i_n228 = axilite_i_axilite_bvalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:441:28  */
  assign axilite_i_n229 = axilite_i_axilite_bresp_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:443:24  */
  assign axilite_i_n230 = axilite_i_bus_waddr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:444:24  */
  assign axilite_i_n231 = axilite_i_bus_raddr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:445:24  */
  assign axilite_i_n232 = axilite_i_bus_write_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:446:23  */
  assign axilite_i_n233 = axilite_i_bus_read_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:447:28  */
  assign axilite_i_n234 = axilite_i_bus_writedata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:419:1  */
  axilite axilite_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .axilite_araddr_in(axilite_araddr_in),
    .axilite_arvalid_in(axilite_arvalid_in),
    .axilite_rready_in(axilite_rready_in),
    .axilite_awaddr_in(axilite_awaddr_in),
    .axilite_awvalid_in(axilite_awvalid_in),
    .axilite_wvalid_in(axilite_wvalid_in),
    .axilite_wdata_in(axilite_wdata_in),
    .axilite_bready_in(axilite_bready_in),
    .bus_readdata_in(host_readdata),
    .bus_readdatavalid_in(host_readdatavalid),
    .bus_writewait_in(host_writewait),
    .bus_readwait_in(host_readwait),
    .axilite_arready_out(axilite_i_axilite_arready_out),
    .axilite_rvalid_out(axilite_i_axilite_rvalid_out),
    .axilite_rlast_out(axilite_i_axilite_rlast_out),
    .axilite_rdata_out(axilite_i_axilite_rdata_out),
    .axilite_rresp_out(axilite_i_axilite_rresp_out),
    .axilite_awready_out(axilite_i_axilite_awready_out),
    .axilite_wready_out(axilite_i_axilite_wready_out),
    .axilite_bvalid_out(axilite_i_axilite_bvalid_out),
    .axilite_bresp_out(axilite_i_axilite_bresp_out),
    .bus_waddr_out(axilite_i_bus_waddr_out),
    .bus_raddr_out(axilite_i_bus_raddr_out),
    .bus_write_out(axilite_i_bus_write_out),
    .bus_read_out(axilite_i_bus_read_out),
    .bus_writedata_out(axilite_i_bus_writedata_out));
  /* ../../HW/src/top/ztachip.vhd:474:33  */
  assign sram_i_n263 = sram_i_dp_readdatavalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:475:36  */
  assign sram_i_n264 = sram_i_dp_readdatavalid_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:476:28  */
  assign sram_i_n265 = sram_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:458:1  */
  sram_core sram_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .dp_rd_addr_in(sram_read_addr),
    .dp_wr_addr_in(sram_write_addr),
    .dp_rd_fork_in(sram_read_fork),
    .dp_wr_fork_in(sram_write_fork),
    .dp_write_in(sram_write_enable),
    .dp_write_vector_in(sram_write_vector),
    .dp_read_in(sram_read_enable),
    .dp_read_vm_in(sram_read_vm),
    .dp_read_vector_in(sram_read_vector),
    .dp_read_gen_valid_in(sram_read_gen_valid),
    .dp_writedata_in(sram_write_data),
    .dp_readdatavalid_out(sram_i_dp_readdatavalid_out),
    .dp_readdatavalid_vm_out(sram_i_dp_readdatavalid_vm_out),
    .dp_readdata_out(sram_i_dp_readdata_out));
  /* ../../HW/src/top/ztachip.vhd:485:34  */
  assign n272_o = ddr_read_wait & ddr_read_enable;
  /* ../../HW/src/top/ztachip.vhd:486:71  */
  assign n274_o = ~ddr_read_wait;
  /* ../../HW/src/top/ztachip.vhd:486:53  */
  assign n275_o = n274_o & ddr_read_enable;
  /* ../../HW/src/top/ztachip.vhd:486:26  */
  assign n276_o = n275_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ztachip.vhd:490:36  */
  assign n278_o = ddr_write_wait & ddr_write_enable;
  /* ../../HW/src/top/ztachip.vhd:491:74  */
  assign n280_o = ~ddr_write_wait;
  /* ../../HW/src/top/ztachip.vhd:491:55  */
  assign n281_o = n280_o & ddr_write_enable;
  /* ../../HW/src/top/ztachip.vhd:491:27  */
  assign n282_o = n281_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ztachip.vhd:495:21  */
  assign n286_o = ~ddr_data_ready;
  /* ../../HW/src/top/ztachip.vhd:495:1  */
  assign n289_o = n286_o ? 1'b1 : 1'b0;
  /* ../../HW/src/top/ztachip.vhd:519:30  */
  assign ddr_rx_i_n292 = ddr_rx_i_read_data_ready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:524:30  */
  assign ddr_rx_i_n294 = ddr_rx_i_read_data_valid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:525:33  */
  assign ddr_rx_i_n295 = ddr_rx_i_read_data_valid_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:526:24  */
  assign ddr_rx_i_n296 = ddr_rx_i_read_data_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:527:32  */
  assign ddr_rx_i_n297 = ddr_rx_i_read_wait_request_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:530:25  */
  assign ddr_rx_i_n298 = ddr_rx_i_ddr_araddr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:531:24  */
  assign ddr_rx_i_n299 = ddr_rx_i_ddr_arlen_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:532:26  */
  assign ddr_rx_i_n300 = ddr_rx_i_ddr_arvalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:537:25  */
  assign ddr_rx_i_n301 = ddr_rx_i_ddr_rready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:538:26  */
  assign ddr_rx_i_n302 = ddr_rx_i_ddr_arburst_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:539:26  */
  assign ddr_rx_i_n303 = ddr_rx_i_ddr_arcache_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:540:23  */
  assign ddr_rx_i_n304 = ddr_rx_i_ddr_arid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:541:25  */
  assign ddr_rx_i_n305 = ddr_rx_i_ddr_arlock_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:542:25  */
  assign ddr_rx_i_n306 = ddr_rx_i_ddr_arprot_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:543:24  */
  assign ddr_rx_i_n307 = ddr_rx_i_ddr_arqos_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:544:25  */
  assign ddr_rx_i_n308 = ddr_rx_i_ddr_arsize_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:506:1  */
  ddr_rx ddr_rx_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .read_addr_in(ddr_read_addr),
    .read_cs_in(ddr_read_enable_2),
    .read_in(ddr_read_enable_2),
    .read_vm_in(ddr_read_vm),
    .read_vector_in(ddr_read_vector),
    .read_fork_in(n291_o),
    .read_start_in(ddr_read_start),
    .read_end_in(ddr_read_end),
    .read_data_wait_in(ddr_data_wait),
    .read_burstlen_in(ddr_read_burstlen),
    .read_filler_data_in(ddr_read_filler_data),
    .ddr_rvalid_in(axi_rvalid_in),
    .ddr_rlast_in(axi_rlast_in),
    .ddr_rdata_in(axi_rdata_in),
    .ddr_arready_in(axi_arready_in),
    .read_data_ready_out(ddr_rx_i_read_data_ready_out),
    .read_fork_out(),
    .read_data_valid_out(ddr_rx_i_read_data_valid_out),
    .read_data_valid_vm_out(ddr_rx_i_read_data_valid_vm_out),
    .read_data_out(ddr_rx_i_read_data_out),
    .read_wait_request_out(ddr_rx_i_read_wait_request_out),
    .ddr_araddr_out(ddr_rx_i_ddr_araddr_out),
    .ddr_arlen_out(ddr_rx_i_ddr_arlen_out),
    .ddr_arvalid_out(ddr_rx_i_ddr_arvalid_out),
    .ddr_rready_out(ddr_rx_i_ddr_rready_out),
    .ddr_arburst_out(ddr_rx_i_ddr_arburst_out),
    .ddr_arcache_out(ddr_rx_i_ddr_arcache_out),
    .ddr_arid_out(ddr_rx_i_ddr_arid_out),
    .ddr_arlock_out(ddr_rx_i_ddr_arlock_out),
    .ddr_arprot_out(ddr_rx_i_ddr_arprot_out),
    .ddr_arqos_out(ddr_rx_i_ddr_arqos_out),
    .ddr_arsize_out(ddr_rx_i_ddr_arsize_out));
  /* ../../HW/src/top/ztachip.vhd:562:33  */
  assign ddr_tx_i_n342 = ddr_tx_i_write_wait_request_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:567:25  */
  assign ddr_tx_i_n343 = ddr_tx_i_ddr_awaddr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:568:24  */
  assign ddr_tx_i_n344 = ddr_tx_i_ddr_awlen_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:569:26  */
  assign ddr_tx_i_n345 = ddr_tx_i_ddr_awvalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:570:24  */
  assign ddr_tx_i_n346 = ddr_tx_i_ddr_waddr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:571:25  */
  assign ddr_tx_i_n347 = ddr_tx_i_ddr_wvalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:572:24  */
  assign ddr_tx_i_n348 = ddr_tx_i_ddr_wdata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:573:24  */
  assign ddr_tx_i_n349 = ddr_tx_i_ddr_wlast_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:574:22  */
  assign ddr_tx_i_n350 = ddr_tx_i_ddr_wbe_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:578:26  */
  assign ddr_tx_i_n351 = ddr_tx_i_ddr_awburst_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:579:26  */
  assign ddr_tx_i_n352 = ddr_tx_i_ddr_awcache_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:580:23  */
  assign ddr_tx_i_n353 = ddr_tx_i_ddr_awid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:581:25  */
  assign ddr_tx_i_n354 = ddr_tx_i_ddr_awlock_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:582:25  */
  assign ddr_tx_i_n355 = ddr_tx_i_ddr_awprot_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:583:24  */
  assign ddr_tx_i_n356 = ddr_tx_i_ddr_awqos_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:584:25  */
  assign ddr_tx_i_n357 = ddr_tx_i_ddr_awsize_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:585:25  */
  assign ddr_tx_i_n358 = ddr_tx_i_ddr_bready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:587:26  */
  assign ddr_tx_i_n359 = ddr_tx_i_ddr_tx_busy_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:551:1  */
  ddr_tx ddr_tx_i (
    .clock_in(clock_in),
    .reset_in(reset_in),
    .write_addr_in(ddr_write_addr),
    .write_cs_in(ddr_write_enable_2),
    .write_in(ddr_write_enable_2),
    .write_vector_in(ddr_write_vector),
    .write_end_in(ddr_write_end),
    .write_data_in(ddr_write_data),
    .write_burstlen_in(ddr_write_burstlen),
    .write_burstlen2_in(ddr_write_burstlen2),
    .write_burstlen3_in(ddr_write_burstlen3),
    .ddr_awready_in(axi_awready_in),
    .ddr_wready_in(axi_wready_in),
    .ddr_bresp_in(axi_bresp_in),
    .write_wait_request_out(ddr_tx_i_write_wait_request_out),
    .ddr_awaddr_out(ddr_tx_i_ddr_awaddr_out),
    .ddr_awlen_out(ddr_tx_i_ddr_awlen_out),
    .ddr_awvalid_out(ddr_tx_i_ddr_awvalid_out),
    .ddr_waddr_out(ddr_tx_i_ddr_waddr_out),
    .ddr_wvalid_out(ddr_tx_i_ddr_wvalid_out),
    .ddr_wdata_out(ddr_tx_i_ddr_wdata_out),
    .ddr_wlast_out(ddr_tx_i_ddr_wlast_out),
    .ddr_wbe_out(ddr_tx_i_ddr_wbe_out),
    .ddr_awburst_out(ddr_tx_i_ddr_awburst_out),
    .ddr_awcache_out(ddr_tx_i_ddr_awcache_out),
    .ddr_awid_out(ddr_tx_i_ddr_awid_out),
    .ddr_awlock_out(ddr_tx_i_ddr_awlock_out),
    .ddr_awprot_out(ddr_tx_i_ddr_awprot_out),
    .ddr_awqos_out(ddr_tx_i_ddr_awqos_out),
    .ddr_awsize_out(ddr_tx_i_ddr_awsize_out),
    .ddr_bready_out(ddr_tx_i_ddr_bready_out),
    .ddr_tx_busy_out(ddr_tx_i_ddr_tx_busy_out));
  /* ../../HW/src/top/ztachip.vhd:603:33  */
  assign n396_o = host_waddr[13:2];
  /* ../../HW/src/top/ztachip.vhd:604:33  */
  assign n397_o = host_raddr[13:2];
  /* ../../HW/src/top/ztachip.vhd:608:27  */
  assign dp_1_i_n398 = dp_1_i_bus_readdata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:609:32  */
  assign dp_1_i_n399 = dp_1_i_bus_readdatavalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:610:28  */
  assign dp_1_i_n400 = dp_1_i_bus_writewait_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:611:27  */
  assign dp_1_i_n401 = dp_1_i_bus_readwait_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:615:31  */
  assign dp_1_i_n402 = dp_1_i_readmaster1_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:616:31  */
  assign dp_1_i_n403 = dp_1_i_readmaster1_fork_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:617:36  */
  assign dp_1_i_n404 = dp_1_i_readmaster1_addr_mode_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:619:31  */
  assign dp_1_i_n406 = dp_1_i_readmaster1_read_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:620:34  */
  assign dp_1_i_n407 = dp_1_i_readmaster1_read_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:621:41  */
  assign dp_1_i_n408 = dp_1_i_readmaster1_read_data_flow_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:622:38  */
  assign dp_1_i_n409 = dp_1_i_readmaster1_read_stream_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:623:41  */
  assign dp_1_i_n410 = dp_1_i_readmaster1_read_stream_id_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:624:38  */
  assign dp_1_i_n411 = dp_1_i_readmaster1_read_vector_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:625:39  */
  assign dp_1_i_n412 = dp_1_i_readmaster1_read_scatter_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:632:36  */
  assign dp_1_i_n415 = dp_1_i_readmaster1_data_type_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:633:37  */
  assign dp_1_i_n416 = dp_1_i_readmaster1_data_model_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:636:32  */
  assign dp_1_i_n417 = dp_1_i_writemaster1_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:637:32  */
  assign dp_1_i_n418 = dp_1_i_writemaster1_fork_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:638:37  */
  assign dp_1_i_n419 = dp_1_i_writemaster1_addr_mode_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:639:30  */
  assign dp_1_i_n420 = dp_1_i_writemaster1_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:640:33  */
  assign dp_1_i_n421 = dp_1_i_writemaster1_mcast_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:642:33  */
  assign dp_1_i_n423 = dp_1_i_writemaster1_write_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:643:43  */
  assign dp_1_i_n424 = dp_1_i_writemaster1_write_data_flow_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:644:40  */
  assign dp_1_i_n425 = dp_1_i_writemaster1_write_vector_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:645:40  */
  assign dp_1_i_n426 = dp_1_i_writemaster1_write_stream_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:646:43  */
  assign dp_1_i_n427 = dp_1_i_writemaster1_write_stream_id_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:647:41  */
  assign dp_1_i_n428 = dp_1_i_writemaster1_write_scatter_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:648:37  */
  assign dp_1_i_n429 = dp_1_i_writemaster1_writedata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:652:37  */
  assign dp_1_i_n432 = dp_1_i_writemaster1_data_type_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:653:38  */
  assign dp_1_i_n433 = dp_1_i_writemaster1_data_model_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:658:31  */
  assign dp_1_i_n435 = dp_1_i_readmaster2_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:659:31  */
  assign dp_1_i_n436 = dp_1_i_readmaster2_fork_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:661:31  */
  assign dp_1_i_n438 = dp_1_i_readmaster2_read_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:662:34  */
  assign dp_1_i_n439 = dp_1_i_readmaster2_read_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:663:38  */
  assign dp_1_i_n440 = dp_1_i_readmaster2_read_vector_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:674:32  */
  assign dp_1_i_n444 = dp_1_i_writemaster2_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:675:32  */
  assign dp_1_i_n445 = dp_1_i_writemaster2_fork_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:677:33  */
  assign dp_1_i_n447 = dp_1_i_writemaster2_write_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:678:30  */
  assign dp_1_i_n448 = dp_1_i_writemaster2_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:679:40  */
  assign dp_1_i_n449 = dp_1_i_writemaster2_write_vector_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:681:37  */
  assign dp_1_i_n451 = dp_1_i_writemaster2_writedata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:690:31  */
  assign dp_1_i_n455 = dp_1_i_readmaster3_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:692:31  */
  assign dp_1_i_n457 = dp_1_i_readmaster3_read_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:693:34  */
  assign dp_1_i_n458 = dp_1_i_readmaster3_read_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:694:38  */
  assign dp_1_i_n459 = dp_1_i_readmaster3_read_vector_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:696:37  */
  assign dp_1_i_n461 = dp_1_i_readmaster3_read_start_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:697:35  */
  assign dp_1_i_n462 = dp_1_i_readmaster3_read_end_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:702:35  */
  assign dp_1_i_n463 = dp_1_i_readmaster3_burstlen_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:704:38  */
  assign dp_1_i_n465 = dp_1_i_readmaster3_filler_data_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:707:32  */
  assign dp_1_i_n466 = dp_1_i_writemaster3_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:709:33  */
  assign dp_1_i_n468 = dp_1_i_writemaster3_write_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:711:40  */
  assign dp_1_i_n470 = dp_1_i_writemaster3_write_vector_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:713:37  */
  assign dp_1_i_n472 = dp_1_i_writemaster3_write_end_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:714:37  */
  assign dp_1_i_n473 = dp_1_i_writemaster3_writedata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:716:36  */
  assign dp_1_i_n474 = dp_1_i_writemaster3_burstlen_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:717:37  */
  assign dp_1_i_n475 = dp_1_i_writemaster3_burstlen2_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:718:37  */
  assign dp_1_i_n476 = dp_1_i_writemaster3_burstlen3_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:724:30  */
  assign dp_1_i_n479 = dp_1_i_task_start_addr_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:725:19  */
  assign dp_1_i_n480 = dp_1_i_task_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:726:22  */
  assign dp_1_i_n481 = dp_1_i_task_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:727:25  */
  assign dp_1_i_n482 = dp_1_i_task_pcore_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:728:28  */
  assign dp_1_i_n483 = dp_1_i_task_lockstep_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:729:28  */
  assign dp_1_i_n484 = dp_1_i_task_tid_mask_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:730:34  */
  assign dp_1_i_n485 = dp_1_i_task_iregister_auto_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:731:30  */
  assign dp_1_i_n486 = dp_1_i_task_data_model_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:734:24  */
  assign dp_1_i_n487 = dp_1_i_task_busy_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:595:1  */
  dp_core dp_1_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .bus_waddr_in(n396_o),
    .bus_raddr_in(n397_o),
    .bus_write_in(host_wren),
    .bus_read_in(host_rden),
    .bus_writedata_in(host_writedata),
    .readmaster1_readdatavalid_in(pcore_read_data_valid2),
    .readmaster1_readdatavalid_vm_in(pcore_readdata_vm),
    .readmaster1_readdata_in(pcore_read_data),
    .readmaster1_wait_request_in(dp_pcore_read_wait),
    .writemaster1_wait_request_in(dp_pcore_write_wait),
    .writemaster1_counter_in(pcore_write_counter_r),
    .readmaster2_readdatavalid_in(sram_read_data_valid),
    .readmaster2_readdatavalid_vm_in(sram_readdata_vm),
    .readmaster2_readdata_in(sram_read_data),
    .readmaster2_wait_request_in(dp_sram_read_wait),
    .writemaster2_wait_request_in(dp_sram_write_wait),
    .writemaster2_counter_in(sram_write_counter_r),
    .readmaster3_readdatavalid_in(ddr_read_data_valid),
    .readmaster3_readdatavalid_vm_in(ddr_readdata_vm),
    .readmaster3_readdata_in(ddr_read_data),
    .readmaster3_wait_request_in(ddr_read_wait_2),
    .writemaster3_wait_request_in(ddr_write_wait_2),
    .writemaster3_counter_in(ddr_write_counter_r),
    .task_busy_in(busy),
    .task_ready_in(ready),
    .bar_in(bar),
    .ddr_tx_busy_in(ddr_tx_busy),
    .bus_readdata_out(dp_1_i_bus_readdata_out),
    .bus_readdatavalid_out(dp_1_i_bus_readdatavalid_out),
    .bus_writewait_out(dp_1_i_bus_writewait_out),
    .bus_readwait_out(dp_1_i_bus_readwait_out),
    .readmaster1_addr_out(dp_1_i_readmaster1_addr_out),
    .readmaster1_fork_out(dp_1_i_readmaster1_fork_out),
    .readmaster1_addr_mode_out(dp_1_i_readmaster1_addr_mode_out),
    .readmaster1_cs_out(),
    .readmaster1_read_out(dp_1_i_readmaster1_read_out),
    .readmaster1_read_vm_out(dp_1_i_readmaster1_read_vm_out),
    .readmaster1_read_data_flow_out(dp_1_i_readmaster1_read_data_flow_out),
    .readmaster1_read_stream_out(dp_1_i_readmaster1_read_stream_out),
    .readmaster1_read_stream_id_out(dp_1_i_readmaster1_read_stream_id_out),
    .readmaster1_read_vector_out(dp_1_i_readmaster1_read_vector_out),
    .readmaster1_read_scatter_out(dp_1_i_readmaster1_read_scatter_out),
    .readmaster1_burstlen_out(),
    .readmaster1_bus_id_out(),
    .readmaster1_data_type_out(dp_1_i_readmaster1_data_type_out),
    .readmaster1_data_model_out(dp_1_i_readmaster1_data_model_out),
    .writemaster1_addr_out(dp_1_i_writemaster1_addr_out),
    .writemaster1_fork_out(dp_1_i_writemaster1_fork_out),
    .writemaster1_addr_mode_out(dp_1_i_writemaster1_addr_mode_out),
    .writemaster1_vm_out(dp_1_i_writemaster1_vm_out),
    .writemaster1_mcast_out(dp_1_i_writemaster1_mcast_out),
    .writemaster1_cs_out(),
    .writemaster1_write_out(dp_1_i_writemaster1_write_out),
    .writemaster1_write_data_flow_out(dp_1_i_writemaster1_write_data_flow_out),
    .writemaster1_write_vector_out(dp_1_i_writemaster1_write_vector_out),
    .writemaster1_write_stream_out(dp_1_i_writemaster1_write_stream_out),
    .writemaster1_write_stream_id_out(dp_1_i_writemaster1_write_stream_id_out),
    .writemaster1_write_scatter_out(dp_1_i_writemaster1_write_scatter_out),
    .writemaster1_writedata_out(dp_1_i_writemaster1_writedata_out),
    .writemaster1_burstlen_out(),
    .writemaster1_bus_id_out(),
    .writemaster1_data_type_out(dp_1_i_writemaster1_data_type_out),
    .writemaster1_data_model_out(dp_1_i_writemaster1_data_model_out),
    .writemaster1_thread_out(),
    .readmaster2_addr_out(dp_1_i_readmaster2_addr_out),
    .readmaster2_fork_out(dp_1_i_readmaster2_fork_out),
    .readmaster2_cs_out(),
    .readmaster2_read_out(dp_1_i_readmaster2_read_out),
    .readmaster2_read_vm_out(dp_1_i_readmaster2_read_vm_out),
    .readmaster2_read_vector_out(dp_1_i_readmaster2_read_vector_out),
    .readmaster2_read_scatter_out(),
    .readmaster2_burstlen_out(),
    .readmaster2_bus_id_out(),
    .writemaster2_addr_out(dp_1_i_writemaster2_addr_out),
    .writemaster2_fork_out(dp_1_i_writemaster2_fork_out),
    .writemaster2_cs_out(),
    .writemaster2_write_out(dp_1_i_writemaster2_write_out),
    .writemaster2_vm_out(dp_1_i_writemaster2_vm_out),
    .writemaster2_write_vector_out(dp_1_i_writemaster2_write_vector_out),
    .writemaster2_write_scatter_out(),
    .writemaster2_writedata_out(dp_1_i_writemaster2_writedata_out),
    .writemaster2_burstlen_out(),
    .writemaster2_bus_id_out(),
    .writemaster2_thread_out(),
    .readmaster3_addr_out(dp_1_i_readmaster3_addr_out),
    .readmaster3_cs_out(),
    .readmaster3_read_out(dp_1_i_readmaster3_read_out),
    .readmaster3_read_vm_out(dp_1_i_readmaster3_read_vm_out),
    .readmaster3_read_vector_out(dp_1_i_readmaster3_read_vector_out),
    .readmaster3_read_scatter_out(),
    .readmaster3_read_start_out(dp_1_i_readmaster3_read_start_out),
    .readmaster3_read_end_out(dp_1_i_readmaster3_read_end_out),
    .readmaster3_burstlen_out(dp_1_i_readmaster3_burstlen_out),
    .readmaster3_bus_id_out(),
    .readmaster3_filler_data_out(dp_1_i_readmaster3_filler_data_out),
    .writemaster3_addr_out(dp_1_i_writemaster3_addr_out),
    .writemaster3_cs_out(),
    .writemaster3_write_out(dp_1_i_writemaster3_write_out),
    .writemaster3_vm_out(),
    .writemaster3_write_vector_out(dp_1_i_writemaster3_write_vector_out),
    .writemaster3_write_scatter_out(),
    .writemaster3_write_end_out(dp_1_i_writemaster3_write_end_out),
    .writemaster3_writedata_out(dp_1_i_writemaster3_writedata_out),
    .writemaster3_burstlen_out(dp_1_i_writemaster3_burstlen_out),
    .writemaster3_burstlen2_out(dp_1_i_writemaster3_burstlen2_out),
    .writemaster3_burstlen3_out(dp_1_i_writemaster3_burstlen3_out),
    .writemaster3_bus_id_out(),
    .writemaster3_thread_out(),
    .writemaster3_filler_data_out(),
    .task_start_addr_out(dp_1_i_task_start_addr_out),
    .task_out(dp_1_i_task_out),
    .task_vm_out(dp_1_i_task_vm_out),
    .task_pcore_out(dp_1_i_task_pcore_out),
    .task_lockstep_out(dp_1_i_task_lockstep_out),
    .task_tid_mask_out(dp_1_i_task_tid_mask_out),
    .task_iregister_auto_out(dp_1_i_task_iregister_auto_out),
    .task_data_model_out(dp_1_i_task_data_model_out),
    .task_busy_out(dp_1_i_task_busy_out),
    .indication_avail_out());
  /* ../../HW/src/top/ztachip.vhd:766:30  */
  assign core_i_n646 = core_i_dp_write_wait_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:777:29  */
  assign core_i_n647 = core_i_dp_read_wait_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:786:32  */
  assign core_i_n648 = core_i_dp_readdatavalid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:787:33  */
  assign core_i_n649 = core_i_dp_read_gen_valid_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:788:28  */
  assign core_i_n650 = core_i_dp_readdata_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:789:29  */
  assign core_i_n651 = core_i_dp_readdata_vm_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:802:21  */
  assign core_i_n652 = core_i_busy_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:803:22  */
  assign core_i_n653 = core_i_ready_out; // (signal)
  /* ../../HW/src/top/ztachip.vhd:750:1  */
  core core_i (
    .clock_in(clock_in),
    .clock_x2_in(clock_x2_in),
    .reset_in(reset_in),
    .dp_rd_addr_in(pcore_read_addr),
    .dp_rd_fork_in(pcore_read_fork),
    .dp_rd_addr_mode_in(pcore_read_addr_mode),
    .dp_wr_addr_in(pcore_write_addr),
    .dp_wr_fork_in(pcore_write_fork),
    .dp_wr_addr_mode_in(pcore_write_addr_mode),
    .dp_wr_mcast_in(pcore_mcast),
    .dp_write_in(pcore_write_enable),
    .dp_write_data_flow_in(pcore_write_data_flow),
    .dp_write_data_type_in(pcore_write_data_type),
    .dp_write_data_model_in(pcore_write_data_model),
    .dp_write_gen_valid_in(pcore_write_gen_valid),
    .dp_write_vector_in(pcore_write_vector),
    .dp_write_stream_in(pcore_write_stream),
    .dp_write_stream_id_in(pcore_write_stream_id),
    .dp_write_scatter_in(pcore_write_scatter2),
    .dp_read_gen_valid_in(pcore_read_gen_valid),
    .dp_read_in(pcore_read_enable),
    .dp_read_data_flow_in(pcore_read_data_flow),
    .dp_read_stream_in(pcore_read_stream),
    .dp_read_stream_id_in(pcore_read_stream_id),
    .dp_read_data_type_in(pcore_read_data_type),
    .dp_read_data_model_in(pcore_read_data_model),
    .dp_read_vector_in(pcore_read_vector),
    .dp_read_scatter_in(pcore_read_scatter2),
    .dp_writedata_in(pcore_write_data),
    .task_start_addr_in(task_start_addr),
    .task_in(\task ),
    .task_vm_in(task_vm),
    .task_pcore_in(task_pcore),
    .task_lockstep_in(task_lockstep),
    .task_tid_mask_in(task_tid_mask),
    .task_iregister_auto_in(task_iregister_auto),
    .task_data_model_in(task_data_model),
    .dp_write_wait_out(core_i_dp_write_wait_out),
    .dp_read_wait_out(core_i_dp_read_wait_out),
    .dp_readdatavalid_out(core_i_dp_readdatavalid_out),
    .dp_read_gen_valid_out(core_i_dp_read_gen_valid_out),
    .dp_readdata_out(core_i_dp_readdata_out),
    .dp_readdata_vm_out(core_i_dp_readdata_vm_out),
    .busy_out(core_i_busy_out),
    .ready_out(core_i_ready_out));
  assign n670_o = {1'b0, 23'b00000000000000000000000, 24'b000000000000000000000000, 24'b000000000000000000000000};
  /* ../../HW/src/top/ztachip.vhd:367:9  */
  assign n671_o = n82_o ? n127_o : pcore_write_counter_r;
  /* ../../HW/src/top/ztachip.vhd:367:9  */
  always @(posedge clock_in or posedge n79_o)
    if (n79_o)
      n672_q <= 48'b000000000000000000000000000000000000000000000000;
    else
      n672_q <= n671_o;
  /* ../../HW/src/top/ztachip.vhd:367:9  */
  assign n673_o = n131_o ? n176_o : sram_write_counter_r;
  /* ../../HW/src/top/ztachip.vhd:367:9  */
  always @(posedge clock_in or posedge n79_o)
    if (n79_o)
      n674_q <= 48'b000000000000000000000000000000000000000000000000;
    else
      n674_q <= n673_o;
  /* ../../HW/src/top/ztachip.vhd:367:9  */
  assign n675_o = n180_o ? n197_o : ddr_write_counter_r;
  /* ../../HW/src/top/ztachip.vhd:367:9  */
  always @(posedge clock_in or posedge n79_o)
    if (n79_o)
      n676_q <= 24'b000000000000000000000000;
    else
      n676_q <= n675_o;
  /* ../../HW/src/top/ztachip.vhd:803:22  */
  assign n678_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:802:21  */
  assign n679_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:375:72  */
  assign n680_o = n91_o ? n679_o : n678_o;
  /* ../../HW/src/top/ztachip.vhd:375:20  */
  assign n681_o = n89_o;
  /* ../../HW/src/top/ztachip.vhd:375:20  */
  assign n682_o = ~n681_o;
  /* ../../HW/src/top/ztachip.vhd:788:28  */
  assign n683_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:375:20  */
  assign n684_o = n682_o ? n95_o : n683_o;
  /* ../../HW/src/top/ztachip.vhd:786:32  */
  assign n685_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:375:20  */
  assign n686_o = n681_o ? n95_o : n685_o;
  /* ../../HW/src/top/ztachip.vhd:766:30  */
  assign n687_o = {n686_o, n684_o};
  /* ../../HW/src/top/ztachip.vhd:375:42  */
  assign n688_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:375:20  */
  assign n689_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:377:72  */
  assign n690_o = n101_o ? n689_o : n688_o;
  /* ../../HW/src/top/ztachip.vhd:377:20  */
  assign n691_o = n99_o;
  /* ../../HW/src/top/ztachip.vhd:377:20  */
  assign n692_o = ~n691_o;
  /* ../../HW/src/top/ztachip.vhd:750:1  */
  assign n693_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:377:20  */
  assign n694_o = n692_o ? n105_o : n693_o;
  /* ../../HW/src/top/ztachip.vhd:750:1  */
  assign n695_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:377:20  */
  assign n696_o = n691_o ? n105_o : n695_o;
  /* ../../HW/src/top/ztachip.vhd:750:1  */
  assign n697_o = {n696_o, n694_o};
  /* ../../HW/src/top/ztachip.vhd:377:42  */
  assign n698_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:377:20  */
  assign n699_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:379:72  */
  assign n700_o = n111_o ? n699_o : n698_o;
  /* ../../HW/src/top/ztachip.vhd:379:20  */
  assign n701_o = n109_o;
  /* ../../HW/src/top/ztachip.vhd:379:20  */
  assign n702_o = ~n701_o;
  /* ../../HW/src/top/ztachip.vhd:750:1  */
  assign n703_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:379:20  */
  assign n704_o = n702_o ? n115_o : n703_o;
  /* ../../HW/src/top/ztachip.vhd:731:30  */
  assign n705_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:379:20  */
  assign n706_o = n701_o ? n115_o : n705_o;
  /* ../../HW/src/top/ztachip.vhd:729:28  */
  assign n707_o = {n706_o, n704_o};
  /* ../../HW/src/top/ztachip.vhd:379:42  */
  assign n708_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:379:20  */
  assign n709_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:381:72  */
  assign n710_o = n119_o ? n709_o : n708_o;
  /* ../../HW/src/top/ztachip.vhd:381:20  */
  assign n711_o = n117_o;
  /* ../../HW/src/top/ztachip.vhd:381:20  */
  assign n712_o = ~n711_o;
  /* ../../HW/src/top/ztachip.vhd:727:25  */
  assign n713_o = pcore_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:381:20  */
  assign n714_o = n712_o ? n123_o : n713_o;
  /* ../../HW/src/top/ztachip.vhd:725:19  */
  assign n715_o = pcore_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:381:20  */
  assign n716_o = n711_o ? n123_o : n715_o;
  /* ../../HW/src/top/ztachip.vhd:718:37  */
  assign n717_o = {n716_o, n714_o};
  /* ../../HW/src/top/ztachip.vhd:381:42  */
  assign n718_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:381:20  */
  assign n719_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:391:75  */
  assign n720_o = n140_o ? n719_o : n718_o;
  /* ../../HW/src/top/ztachip.vhd:391:20  */
  assign n721_o = n138_o;
  /* ../../HW/src/top/ztachip.vhd:391:20  */
  assign n722_o = ~n721_o;
  /* ../../HW/src/top/ztachip.vhd:716:36  */
  assign n723_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:391:20  */
  assign n724_o = n722_o ? n144_o : n723_o;
  /* ../../HW/src/top/ztachip.vhd:713:37  */
  assign n725_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:391:20  */
  assign n726_o = n721_o ? n144_o : n725_o;
  /* ../../HW/src/top/ztachip.vhd:709:33  */
  assign n727_o = {n726_o, n724_o};
  /* ../../HW/src/top/ztachip.vhd:391:41  */
  assign n728_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:391:20  */
  assign n729_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:393:75  */
  assign n730_o = n150_o ? n729_o : n728_o;
  /* ../../HW/src/top/ztachip.vhd:393:20  */
  assign n731_o = n148_o;
  /* ../../HW/src/top/ztachip.vhd:393:20  */
  assign n732_o = ~n731_o;
  /* ../../HW/src/top/ztachip.vhd:704:38  */
  assign n733_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:393:20  */
  assign n734_o = n732_o ? n154_o : n733_o;
  /* ../../HW/src/top/ztachip.vhd:697:35  */
  assign n735_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:393:20  */
  assign n736_o = n731_o ? n154_o : n735_o;
  /* ../../HW/src/top/ztachip.vhd:694:38  */
  assign n737_o = {n736_o, n734_o};
  /* ../../HW/src/top/ztachip.vhd:393:41  */
  assign n738_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:393:20  */
  assign n739_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:395:75  */
  assign n740_o = n160_o ? n739_o : n738_o;
  /* ../../HW/src/top/ztachip.vhd:395:20  */
  assign n741_o = n158_o;
  /* ../../HW/src/top/ztachip.vhd:395:20  */
  assign n742_o = ~n741_o;
  /* ../../HW/src/top/ztachip.vhd:692:31  */
  assign n743_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:395:20  */
  assign n744_o = n742_o ? n164_o : n743_o;
  /* ../../HW/src/top/ztachip.vhd:681:37  */
  assign n745_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:395:20  */
  assign n746_o = n741_o ? n164_o : n745_o;
  /* ../../HW/src/top/ztachip.vhd:678:30  */
  assign n747_o = {n746_o, n744_o};
  /* ../../HW/src/top/ztachip.vhd:395:41  */
  assign n748_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:395:20  */
  assign n749_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:397:75  */
  assign n750_o = n168_o ? n749_o : n748_o;
  /* ../../HW/src/top/ztachip.vhd:397:20  */
  assign n751_o = n166_o;
  /* ../../HW/src/top/ztachip.vhd:397:20  */
  assign n752_o = ~n751_o;
  /* ../../HW/src/top/ztachip.vhd:675:32  */
  assign n753_o = sram_write_counter_r[23:0];
  /* ../../HW/src/top/ztachip.vhd:397:20  */
  assign n754_o = n752_o ? n172_o : n753_o;
  /* ../../HW/src/top/ztachip.vhd:663:38  */
  assign n755_o = sram_write_counter_r[47:24];
  /* ../../HW/src/top/ztachip.vhd:397:20  */
  assign n756_o = n751_o ? n172_o : n755_o;
  /* ../../HW/src/top/ztachip.vhd:661:31  */
  assign n757_o = {n756_o, n754_o};
endmodule

